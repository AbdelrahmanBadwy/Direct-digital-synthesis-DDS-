library ieee;
use ieee.std_logic_1164.all;
-- use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;



entity LUT_DDFS is
	port (
		LUT_line : in  std_logic_vector(15 downto 0);
		LUT_data : out std_logic_vector(15 downto 0) 
	);
end LUT_DDFS;

architecture rtl of LUT_DDFS is
	type LUT_t is array (natural range 0 to 65535) of integer;
	constant LUT: LUT_t := (
		0	=>	32768,
		1	=>	32771,
		2	=>	32774,
		3	=>	32777,
		4	=>	32780,
		5	=>	32783,
		6	=>	32786,
		7	=>	32789,
		8	=>	32793,
		9	=>	32796,
		10	=>	32799,
		11	=>	32802,
		12	=>	32805,
		13	=>	32808,
		14	=>	32811,
		15	=>	32815,
		16	=>	32818,
		17	=>	32821,
		18	=>	32824,
		19	=>	32827,
		20	=>	32830,
		21	=>	32833,
		22	=>	32837,
		23	=>	32840,
		24	=>	32843,
		25	=>	32846,
		26	=>	32849,
		27	=>	32852,
		28	=>	32855,
		29	=>	32859,
		30	=>	32862,
		31	=>	32865,
		32	=>	32868,
		33	=>	32871,
		34	=>	32874,
		35	=>	32877,
		36	=>	32881,
		37	=>	32884,
		38	=>	32887,
		39	=>	32890,
		40	=>	32893,
		41	=>	32896,
		42	=>	32899,
		43	=>	32903,
		44	=>	32906,
		45	=>	32909,
		46	=>	32912,
		47	=>	32915,
		48	=>	32918,
		49	=>	32921,
		50	=>	32925,
		51	=>	32928,
		52	=>	32931,
		53	=>	32934,
		54	=>	32937,
		55	=>	32940,
		56	=>	32943,
		57	=>	32947,
		58	=>	32950,
		59	=>	32953,
		60	=>	32956,
		61	=>	32959,
		62	=>	32962,
		63	=>	32965,
		64	=>	32969,
		65	=>	32972,
		66	=>	32975,
		67	=>	32978,
		68	=>	32981,
		69	=>	32984,
		70	=>	32987,
		71	=>	32991,
		72	=>	32994,
		73	=>	32997,
		74	=>	33000,
		75	=>	33003,
		76	=>	33006,
		77	=>	33009,
		78	=>	33013,
		79	=>	33016,
		80	=>	33019,
		81	=>	33022,
		82	=>	33025,
		83	=>	33028,
		84	=>	33031,
		85	=>	33035,
		86	=>	33038,
		87	=>	33041,
		88	=>	33044,
		89	=>	33047,
		90	=>	33050,
		91	=>	33053,
		92	=>	33057,
		93	=>	33060,
		94	=>	33063,
		95	=>	33066,
		96	=>	33069,
		97	=>	33072,
		98	=>	33075,
		99	=>	33079,
		100	=>	33082,
		101	=>	33085,
		102	=>	33088,
		103	=>	33091,
		104	=>	33094,
		105	=>	33097,
		106	=>	33100,
		107	=>	33104,
		108	=>	33107,
		109	=>	33110,
		110	=>	33113,
		111	=>	33116,
		112	=>	33119,
		113	=>	33122,
		114	=>	33126,
		115	=>	33129,
		116	=>	33132,
		117	=>	33135,
		118	=>	33138,
		119	=>	33141,
		120	=>	33144,
		121	=>	33148,
		122	=>	33151,
		123	=>	33154,
		124	=>	33157,
		125	=>	33160,
		126	=>	33163,
		127	=>	33166,
		128	=>	33170,
		129	=>	33173,
		130	=>	33176,
		131	=>	33179,
		132	=>	33182,
		133	=>	33185,
		134	=>	33188,
		135	=>	33192,
		136	=>	33195,
		137	=>	33198,
		138	=>	33201,
		139	=>	33204,
		140	=>	33207,
		141	=>	33210,
		142	=>	33214,
		143	=>	33217,
		144	=>	33220,
		145	=>	33223,
		146	=>	33226,
		147	=>	33229,
		148	=>	33232,
		149	=>	33236,
		150	=>	33239,
		151	=>	33242,
		152	=>	33245,
		153	=>	33248,
		154	=>	33251,
		155	=>	33254,
		156	=>	33258,
		157	=>	33261,
		158	=>	33264,
		159	=>	33267,
		160	=>	33270,
		161	=>	33273,
		162	=>	33276,
		163	=>	33280,
		164	=>	33283,
		165	=>	33286,
		166	=>	33289,
		167	=>	33292,
		168	=>	33295,
		169	=>	33298,
		170	=>	33302,
		171	=>	33305,
		172	=>	33308,
		173	=>	33311,
		174	=>	33314,
		175	=>	33317,
		176	=>	33320,
		177	=>	33324,
		178	=>	33327,
		179	=>	33330,
		180	=>	33333,
		181	=>	33336,
		182	=>	33339,
		183	=>	33342,
		184	=>	33346,
		185	=>	33349,
		186	=>	33352,
		187	=>	33355,
		188	=>	33358,
		189	=>	33361,
		190	=>	33364,
		191	=>	33368,
		192	=>	33371,
		193	=>	33374,
		194	=>	33377,
		195	=>	33380,
		196	=>	33383,
		197	=>	33386,
		198	=>	33389,
		199	=>	33393,
		200	=>	33396,
		201	=>	33399,
		202	=>	33402,
		203	=>	33405,
		204	=>	33408,
		205	=>	33411,
		206	=>	33415,
		207	=>	33418,
		208	=>	33421,
		209	=>	33424,
		210	=>	33427,
		211	=>	33430,
		212	=>	33433,
		213	=>	33437,
		214	=>	33440,
		215	=>	33443,
		216	=>	33446,
		217	=>	33449,
		218	=>	33452,
		219	=>	33455,
		220	=>	33459,
		221	=>	33462,
		222	=>	33465,
		223	=>	33468,
		224	=>	33471,
		225	=>	33474,
		226	=>	33477,
		227	=>	33481,
		228	=>	33484,
		229	=>	33487,
		230	=>	33490,
		231	=>	33493,
		232	=>	33496,
		233	=>	33499,
		234	=>	33503,
		235	=>	33506,
		236	=>	33509,
		237	=>	33512,
		238	=>	33515,
		239	=>	33518,
		240	=>	33521,
		241	=>	33525,
		242	=>	33528,
		243	=>	33531,
		244	=>	33534,
		245	=>	33537,
		246	=>	33540,
		247	=>	33543,
		248	=>	33547,
		249	=>	33550,
		250	=>	33553,
		251	=>	33556,
		252	=>	33559,
		253	=>	33562,
		254	=>	33565,
		255	=>	33569,
		256	=>	33572,
		257	=>	33575,
		258	=>	33578,
		259	=>	33581,
		260	=>	33584,
		261	=>	33587,
		262	=>	33590,
		263	=>	33594,
		264	=>	33597,
		265	=>	33600,
		266	=>	33603,
		267	=>	33606,
		268	=>	33609,
		269	=>	33612,
		270	=>	33616,
		271	=>	33619,
		272	=>	33622,
		273	=>	33625,
		274	=>	33628,
		275	=>	33631,
		276	=>	33634,
		277	=>	33638,
		278	=>	33641,
		279	=>	33644,
		280	=>	33647,
		281	=>	33650,
		282	=>	33653,
		283	=>	33656,
		284	=>	33660,
		285	=>	33663,
		286	=>	33666,
		287	=>	33669,
		288	=>	33672,
		289	=>	33675,
		290	=>	33678,
		291	=>	33682,
		292	=>	33685,
		293	=>	33688,
		294	=>	33691,
		295	=>	33694,
		296	=>	33697,
		297	=>	33700,
		298	=>	33704,
		299	=>	33707,
		300	=>	33710,
		301	=>	33713,
		302	=>	33716,
		303	=>	33719,
		304	=>	33722,
		305	=>	33726,
		306	=>	33729,
		307	=>	33732,
		308	=>	33735,
		309	=>	33738,
		310	=>	33741,
		311	=>	33744,
		312	=>	33748,
		313	=>	33751,
		314	=>	33754,
		315	=>	33757,
		316	=>	33760,
		317	=>	33763,
		318	=>	33766,
		319	=>	33769,
		320	=>	33773,
		321	=>	33776,
		322	=>	33779,
		323	=>	33782,
		324	=>	33785,
		325	=>	33788,
		326	=>	33791,
		327	=>	33795,
		328	=>	33798,
		329	=>	33801,
		330	=>	33804,
		331	=>	33807,
		332	=>	33810,
		333	=>	33813,
		334	=>	33817,
		335	=>	33820,
		336	=>	33823,
		337	=>	33826,
		338	=>	33829,
		339	=>	33832,
		340	=>	33835,
		341	=>	33839,
		342	=>	33842,
		343	=>	33845,
		344	=>	33848,
		345	=>	33851,
		346	=>	33854,
		347	=>	33857,
		348	=>	33861,
		349	=>	33864,
		350	=>	33867,
		351	=>	33870,
		352	=>	33873,
		353	=>	33876,
		354	=>	33879,
		355	=>	33883,
		356	=>	33886,
		357	=>	33889,
		358	=>	33892,
		359	=>	33895,
		360	=>	33898,
		361	=>	33901,
		362	=>	33905,
		363	=>	33908,
		364	=>	33911,
		365	=>	33914,
		366	=>	33917,
		367	=>	33920,
		368	=>	33923,
		369	=>	33926,
		370	=>	33930,
		371	=>	33933,
		372	=>	33936,
		373	=>	33939,
		374	=>	33942,
		375	=>	33945,
		376	=>	33948,
		377	=>	33952,
		378	=>	33955,
		379	=>	33958,
		380	=>	33961,
		381	=>	33964,
		382	=>	33967,
		383	=>	33970,
		384	=>	33974,
		385	=>	33977,
		386	=>	33980,
		387	=>	33983,
		388	=>	33986,
		389	=>	33989,
		390	=>	33992,
		391	=>	33996,
		392	=>	33999,
		393	=>	34002,
		394	=>	34005,
		395	=>	34008,
		396	=>	34011,
		397	=>	34014,
		398	=>	34018,
		399	=>	34021,
		400	=>	34024,
		401	=>	34027,
		402	=>	34030,
		403	=>	34033,
		404	=>	34036,
		405	=>	34040,
		406	=>	34043,
		407	=>	34046,
		408	=>	34049,
		409	=>	34052,
		410	=>	34055,
		411	=>	34058,
		412	=>	34061,
		413	=>	34065,
		414	=>	34068,
		415	=>	34071,
		416	=>	34074,
		417	=>	34077,
		418	=>	34080,
		419	=>	34083,
		420	=>	34087,
		421	=>	34090,
		422	=>	34093,
		423	=>	34096,
		424	=>	34099,
		425	=>	34102,
		426	=>	34105,
		427	=>	34109,
		428	=>	34112,
		429	=>	34115,
		430	=>	34118,
		431	=>	34121,
		432	=>	34124,
		433	=>	34127,
		434	=>	34131,
		435	=>	34134,
		436	=>	34137,
		437	=>	34140,
		438	=>	34143,
		439	=>	34146,
		440	=>	34149,
		441	=>	34153,
		442	=>	34156,
		443	=>	34159,
		444	=>	34162,
		445	=>	34165,
		446	=>	34168,
		447	=>	34171,
		448	=>	34174,
		449	=>	34178,
		450	=>	34181,
		451	=>	34184,
		452	=>	34187,
		453	=>	34190,
		454	=>	34193,
		455	=>	34196,
		456	=>	34200,
		457	=>	34203,
		458	=>	34206,
		459	=>	34209,
		460	=>	34212,
		461	=>	34215,
		462	=>	34218,
		463	=>	34222,
		464	=>	34225,
		465	=>	34228,
		466	=>	34231,
		467	=>	34234,
		468	=>	34237,
		469	=>	34240,
		470	=>	34244,
		471	=>	34247,
		472	=>	34250,
		473	=>	34253,
		474	=>	34256,
		475	=>	34259,
		476	=>	34262,
		477	=>	34265,
		478	=>	34269,
		479	=>	34272,
		480	=>	34275,
		481	=>	34278,
		482	=>	34281,
		483	=>	34284,
		484	=>	34287,
		485	=>	34291,
		486	=>	34294,
		487	=>	34297,
		488	=>	34300,
		489	=>	34303,
		490	=>	34306,
		491	=>	34309,
		492	=>	34313,
		493	=>	34316,
		494	=>	34319,
		495	=>	34322,
		496	=>	34325,
		497	=>	34328,
		498	=>	34331,
		499	=>	34335,
		500	=>	34338,
		501	=>	34341,
		502	=>	34344,
		503	=>	34347,
		504	=>	34350,
		505	=>	34353,
		506	=>	34356,
		507	=>	34360,
		508	=>	34363,
		509	=>	34366,
		510	=>	34369,
		511	=>	34372,
		512	=>	34375,
		513	=>	34378,
		514	=>	34382,
		515	=>	34385,
		516	=>	34388,
		517	=>	34391,
		518	=>	34394,
		519	=>	34397,
		520	=>	34400,
		521	=>	34404,
		522	=>	34407,
		523	=>	34410,
		524	=>	34413,
		525	=>	34416,
		526	=>	34419,
		527	=>	34422,
		528	=>	34426,
		529	=>	34429,
		530	=>	34432,
		531	=>	34435,
		532	=>	34438,
		533	=>	34441,
		534	=>	34444,
		535	=>	34447,
		536	=>	34451,
		537	=>	34454,
		538	=>	34457,
		539	=>	34460,
		540	=>	34463,
		541	=>	34466,
		542	=>	34469,
		543	=>	34473,
		544	=>	34476,
		545	=>	34479,
		546	=>	34482,
		547	=>	34485,
		548	=>	34488,
		549	=>	34491,
		550	=>	34495,
		551	=>	34498,
		552	=>	34501,
		553	=>	34504,
		554	=>	34507,
		555	=>	34510,
		556	=>	34513,
		557	=>	34517,
		558	=>	34520,
		559	=>	34523,
		560	=>	34526,
		561	=>	34529,
		562	=>	34532,
		563	=>	34535,
		564	=>	34538,
		565	=>	34542,
		566	=>	34545,
		567	=>	34548,
		568	=>	34551,
		569	=>	34554,
		570	=>	34557,
		571	=>	34560,
		572	=>	34564,
		573	=>	34567,
		574	=>	34570,
		575	=>	34573,
		576	=>	34576,
		577	=>	34579,
		578	=>	34582,
		579	=>	34586,
		580	=>	34589,
		581	=>	34592,
		582	=>	34595,
		583	=>	34598,
		584	=>	34601,
		585	=>	34604,
		586	=>	34607,
		587	=>	34611,
		588	=>	34614,
		589	=>	34617,
		590	=>	34620,
		591	=>	34623,
		592	=>	34626,
		593	=>	34629,
		594	=>	34633,
		595	=>	34636,
		596	=>	34639,
		597	=>	34642,
		598	=>	34645,
		599	=>	34648,
		600	=>	34651,
		601	=>	34655,
		602	=>	34658,
		603	=>	34661,
		604	=>	34664,
		605	=>	34667,
		606	=>	34670,
		607	=>	34673,
		608	=>	34676,
		609	=>	34680,
		610	=>	34683,
		611	=>	34686,
		612	=>	34689,
		613	=>	34692,
		614	=>	34695,
		615	=>	34698,
		616	=>	34702,
		617	=>	34705,
		618	=>	34708,
		619	=>	34711,
		620	=>	34714,
		621	=>	34717,
		622	=>	34720,
		623	=>	34724,
		624	=>	34727,
		625	=>	34730,
		626	=>	34733,
		627	=>	34736,
		628	=>	34739,
		629	=>	34742,
		630	=>	34745,
		631	=>	34749,
		632	=>	34752,
		633	=>	34755,
		634	=>	34758,
		635	=>	34761,
		636	=>	34764,
		637	=>	34767,
		638	=>	34771,
		639	=>	34774,
		640	=>	34777,
		641	=>	34780,
		642	=>	34783,
		643	=>	34786,
		644	=>	34789,
		645	=>	34793,
		646	=>	34796,
		647	=>	34799,
		648	=>	34802,
		649	=>	34805,
		650	=>	34808,
		651	=>	34811,
		652	=>	34814,
		653	=>	34818,
		654	=>	34821,
		655	=>	34824,
		656	=>	34827,
		657	=>	34830,
		658	=>	34833,
		659	=>	34836,
		660	=>	34840,
		661	=>	34843,
		662	=>	34846,
		663	=>	34849,
		664	=>	34852,
		665	=>	34855,
		666	=>	34858,
		667	=>	34861,
		668	=>	34865,
		669	=>	34868,
		670	=>	34871,
		671	=>	34874,
		672	=>	34877,
		673	=>	34880,
		674	=>	34883,
		675	=>	34887,
		676	=>	34890,
		677	=>	34893,
		678	=>	34896,
		679	=>	34899,
		680	=>	34902,
		681	=>	34905,
		682	=>	34909,
		683	=>	34912,
		684	=>	34915,
		685	=>	34918,
		686	=>	34921,
		687	=>	34924,
		688	=>	34927,
		689	=>	34930,
		690	=>	34934,
		691	=>	34937,
		692	=>	34940,
		693	=>	34943,
		694	=>	34946,
		695	=>	34949,
		696	=>	34952,
		697	=>	34956,
		698	=>	34959,
		699	=>	34962,
		700	=>	34965,
		701	=>	34968,
		702	=>	34971,
		703	=>	34974,
		704	=>	34977,
		705	=>	34981,
		706	=>	34984,
		707	=>	34987,
		708	=>	34990,
		709	=>	34993,
		710	=>	34996,
		711	=>	34999,
		712	=>	35003,
		713	=>	35006,
		714	=>	35009,
		715	=>	35012,
		716	=>	35015,
		717	=>	35018,
		718	=>	35021,
		719	=>	35024,
		720	=>	35028,
		721	=>	35031,
		722	=>	35034,
		723	=>	35037,
		724	=>	35040,
		725	=>	35043,
		726	=>	35046,
		727	=>	35050,
		728	=>	35053,
		729	=>	35056,
		730	=>	35059,
		731	=>	35062,
		732	=>	35065,
		733	=>	35068,
		734	=>	35071,
		735	=>	35075,
		736	=>	35078,
		737	=>	35081,
		738	=>	35084,
		739	=>	35087,
		740	=>	35090,
		741	=>	35093,
		742	=>	35097,
		743	=>	35100,
		744	=>	35103,
		745	=>	35106,
		746	=>	35109,
		747	=>	35112,
		748	=>	35115,
		749	=>	35118,
		750	=>	35122,
		751	=>	35125,
		752	=>	35128,
		753	=>	35131,
		754	=>	35134,
		755	=>	35137,
		756	=>	35140,
		757	=>	35144,
		758	=>	35147,
		759	=>	35150,
		760	=>	35153,
		761	=>	35156,
		762	=>	35159,
		763	=>	35162,
		764	=>	35165,
		765	=>	35169,
		766	=>	35172,
		767	=>	35175,
		768	=>	35178,
		769	=>	35181,
		770	=>	35184,
		771	=>	35187,
		772	=>	35191,
		773	=>	35194,
		774	=>	35197,
		775	=>	35200,
		776	=>	35203,
		777	=>	35206,
		778	=>	35209,
		779	=>	35212,
		780	=>	35216,
		781	=>	35219,
		782	=>	35222,
		783	=>	35225,
		784	=>	35228,
		785	=>	35231,
		786	=>	35234,
		787	=>	35238,
		788	=>	35241,
		789	=>	35244,
		790	=>	35247,
		791	=>	35250,
		792	=>	35253,
		793	=>	35256,
		794	=>	35259,
		795	=>	35263,
		796	=>	35266,
		797	=>	35269,
		798	=>	35272,
		799	=>	35275,
		800	=>	35278,
		801	=>	35281,
		802	=>	35285,
		803	=>	35288,
		804	=>	35291,
		805	=>	35294,
		806	=>	35297,
		807	=>	35300,
		808	=>	35303,
		809	=>	35306,
		810	=>	35310,
		811	=>	35313,
		812	=>	35316,
		813	=>	35319,
		814	=>	35322,
		815	=>	35325,
		816	=>	35328,
		817	=>	35332,
		818	=>	35335,
		819	=>	35338,
		820	=>	35341,
		821	=>	35344,
		822	=>	35347,
		823	=>	35350,
		824	=>	35353,
		825	=>	35357,
		826	=>	35360,
		827	=>	35363,
		828	=>	35366,
		829	=>	35369,
		830	=>	35372,
		831	=>	35375,
		832	=>	35378,
		833	=>	35382,
		834	=>	35385,
		835	=>	35388,
		836	=>	35391,
		837	=>	35394,
		838	=>	35397,
		839	=>	35400,
		840	=>	35404,
		841	=>	35407,
		842	=>	35410,
		843	=>	35413,
		844	=>	35416,
		845	=>	35419,
		846	=>	35422,
		847	=>	35425,
		848	=>	35429,
		849	=>	35432,
		850	=>	35435,
		851	=>	35438,
		852	=>	35441,
		853	=>	35444,
		854	=>	35447,
		855	=>	35451,
		856	=>	35454,
		857	=>	35457,
		858	=>	35460,
		859	=>	35463,
		860	=>	35466,
		861	=>	35469,
		862	=>	35472,
		863	=>	35476,
		864	=>	35479,
		865	=>	35482,
		866	=>	35485,
		867	=>	35488,
		868	=>	35491,
		869	=>	35494,
		870	=>	35497,
		871	=>	35501,
		872	=>	35504,
		873	=>	35507,
		874	=>	35510,
		875	=>	35513,
		876	=>	35516,
		877	=>	35519,
		878	=>	35523,
		879	=>	35526,
		880	=>	35529,
		881	=>	35532,
		882	=>	35535,
		883	=>	35538,
		884	=>	35541,
		885	=>	35544,
		886	=>	35548,
		887	=>	35551,
		888	=>	35554,
		889	=>	35557,
		890	=>	35560,
		891	=>	35563,
		892	=>	35566,
		893	=>	35569,
		894	=>	35573,
		895	=>	35576,
		896	=>	35579,
		897	=>	35582,
		898	=>	35585,
		899	=>	35588,
		900	=>	35591,
		901	=>	35595,
		902	=>	35598,
		903	=>	35601,
		904	=>	35604,
		905	=>	35607,
		906	=>	35610,
		907	=>	35613,
		908	=>	35616,
		909	=>	35620,
		910	=>	35623,
		911	=>	35626,
		912	=>	35629,
		913	=>	35632,
		914	=>	35635,
		915	=>	35638,
		916	=>	35641,
		917	=>	35645,
		918	=>	35648,
		919	=>	35651,
		920	=>	35654,
		921	=>	35657,
		922	=>	35660,
		923	=>	35663,
		924	=>	35666,
		925	=>	35670,
		926	=>	35673,
		927	=>	35676,
		928	=>	35679,
		929	=>	35682,
		930	=>	35685,
		931	=>	35688,
		932	=>	35692,
		933	=>	35695,
		934	=>	35698,
		935	=>	35701,
		936	=>	35704,
		937	=>	35707,
		938	=>	35710,
		939	=>	35713,
		940	=>	35717,
		941	=>	35720,
		942	=>	35723,
		943	=>	35726,
		944	=>	35729,
		945	=>	35732,
		946	=>	35735,
		947	=>	35738,
		948	=>	35742,
		949	=>	35745,
		950	=>	35748,
		951	=>	35751,
		952	=>	35754,
		953	=>	35757,
		954	=>	35760,
		955	=>	35763,
		956	=>	35767,
		957	=>	35770,
		958	=>	35773,
		959	=>	35776,
		960	=>	35779,
		961	=>	35782,
		962	=>	35785,
		963	=>	35789,
		964	=>	35792,
		965	=>	35795,
		966	=>	35798,
		967	=>	35801,
		968	=>	35804,
		969	=>	35807,
		970	=>	35810,
		971	=>	35814,
		972	=>	35817,
		973	=>	35820,
		974	=>	35823,
		975	=>	35826,
		976	=>	35829,
		977	=>	35832,
		978	=>	35835,
		979	=>	35839,
		980	=>	35842,
		981	=>	35845,
		982	=>	35848,
		983	=>	35851,
		984	=>	35854,
		985	=>	35857,
		986	=>	35860,
		987	=>	35864,
		988	=>	35867,
		989	=>	35870,
		990	=>	35873,
		991	=>	35876,
		992	=>	35879,
		993	=>	35882,
		994	=>	35885,
		995	=>	35889,
		996	=>	35892,
		997	=>	35895,
		998	=>	35898,
		999	=>	35901,
		1000	=>	35904,
		1001	=>	35907,
		1002	=>	35910,
		1003	=>	35914,
		1004	=>	35917,
		1005	=>	35920,
		1006	=>	35923,
		1007	=>	35926,
		1008	=>	35929,
		1009	=>	35932,
		1010	=>	35936,
		1011	=>	35939,
		1012	=>	35942,
		1013	=>	35945,
		1014	=>	35948,
		1015	=>	35951,
		1016	=>	35954,
		1017	=>	35957,
		1018	=>	35961,
		1019	=>	35964,
		1020	=>	35967,
		1021	=>	35970,
		1022	=>	35973,
		1023	=>	35976,
		1024	=>	35979,
		1025	=>	35982,
		1026	=>	35986,
		1027	=>	35989,
		1028	=>	35992,
		1029	=>	35995,
		1030	=>	35998,
		1031	=>	36001,
		1032	=>	36004,
		1033	=>	36007,
		1034	=>	36011,
		1035	=>	36014,
		1036	=>	36017,
		1037	=>	36020,
		1038	=>	36023,
		1039	=>	36026,
		1040	=>	36029,
		1041	=>	36032,
		1042	=>	36036,
		1043	=>	36039,
		1044	=>	36042,
		1045	=>	36045,
		1046	=>	36048,
		1047	=>	36051,
		1048	=>	36054,
		1049	=>	36057,
		1050	=>	36061,
		1051	=>	36064,
		1052	=>	36067,
		1053	=>	36070,
		1054	=>	36073,
		1055	=>	36076,
		1056	=>	36079,
		1057	=>	36082,
		1058	=>	36086,
		1059	=>	36089,
		1060	=>	36092,
		1061	=>	36095,
		1062	=>	36098,
		1063	=>	36101,
		1064	=>	36104,
		1065	=>	36107,
		1066	=>	36111,
		1067	=>	36114,
		1068	=>	36117,
		1069	=>	36120,
		1070	=>	36123,
		1071	=>	36126,
		1072	=>	36129,
		1073	=>	36132,
		1074	=>	36136,
		1075	=>	36139,
		1076	=>	36142,
		1077	=>	36145,
		1078	=>	36148,
		1079	=>	36151,
		1080	=>	36154,
		1081	=>	36157,
		1082	=>	36161,
		1083	=>	36164,
		1084	=>	36167,
		1085	=>	36170,
		1086	=>	36173,
		1087	=>	36176,
		1088	=>	36179,
		1089	=>	36182,
		1090	=>	36186,
		1091	=>	36189,
		1092	=>	36192,
		1093	=>	36195,
		1094	=>	36198,
		1095	=>	36201,
		1096	=>	36204,
		1097	=>	36207,
		1098	=>	36211,
		1099	=>	36214,
		1100	=>	36217,
		1101	=>	36220,
		1102	=>	36223,
		1103	=>	36226,
		1104	=>	36229,
		1105	=>	36232,
		1106	=>	36236,
		1107	=>	36239,
		1108	=>	36242,
		1109	=>	36245,
		1110	=>	36248,
		1111	=>	36251,
		1112	=>	36254,
		1113	=>	36257,
		1114	=>	36261,
		1115	=>	36264,
		1116	=>	36267,
		1117	=>	36270,
		1118	=>	36273,
		1119	=>	36276,
		1120	=>	36279,
		1121	=>	36282,
		1122	=>	36286,
		1123	=>	36289,
		1124	=>	36292,
		1125	=>	36295,
		1126	=>	36298,
		1127	=>	36301,
		1128	=>	36304,
		1129	=>	36307,
		1130	=>	36311,
		1131	=>	36314,
		1132	=>	36317,
		1133	=>	36320,
		1134	=>	36323,
		1135	=>	36326,
		1136	=>	36329,
		1137	=>	36332,
		1138	=>	36335,
		1139	=>	36339,
		1140	=>	36342,
		1141	=>	36345,
		1142	=>	36348,
		1143	=>	36351,
		1144	=>	36354,
		1145	=>	36357,
		1146	=>	36360,
		1147	=>	36364,
		1148	=>	36367,
		1149	=>	36370,
		1150	=>	36373,
		1151	=>	36376,
		1152	=>	36379,
		1153	=>	36382,
		1154	=>	36385,
		1155	=>	36389,
		1156	=>	36392,
		1157	=>	36395,
		1158	=>	36398,
		1159	=>	36401,
		1160	=>	36404,
		1161	=>	36407,
		1162	=>	36410,
		1163	=>	36414,
		1164	=>	36417,
		1165	=>	36420,
		1166	=>	36423,
		1167	=>	36426,
		1168	=>	36429,
		1169	=>	36432,
		1170	=>	36435,
		1171	=>	36439,
		1172	=>	36442,
		1173	=>	36445,
		1174	=>	36448,
		1175	=>	36451,
		1176	=>	36454,
		1177	=>	36457,
		1178	=>	36460,
		1179	=>	36463,
		1180	=>	36467,
		1181	=>	36470,
		1182	=>	36473,
		1183	=>	36476,
		1184	=>	36479,
		1185	=>	36482,
		1186	=>	36485,
		1187	=>	36488,
		1188	=>	36492,
		1189	=>	36495,
		1190	=>	36498,
		1191	=>	36501,
		1192	=>	36504,
		1193	=>	36507,
		1194	=>	36510,
		1195	=>	36513,
		1196	=>	36517,
		1197	=>	36520,
		1198	=>	36523,
		1199	=>	36526,
		1200	=>	36529,
		1201	=>	36532,
		1202	=>	36535,
		1203	=>	36538,
		1204	=>	36542,
		1205	=>	36545,
		1206	=>	36548,
		1207	=>	36551,
		1208	=>	36554,
		1209	=>	36557,
		1210	=>	36560,
		1211	=>	36563,
		1212	=>	36566,
		1213	=>	36570,
		1214	=>	36573,
		1215	=>	36576,
		1216	=>	36579,
		1217	=>	36582,
		1218	=>	36585,
		1219	=>	36588,
		1220	=>	36591,
		1221	=>	36595,
		1222	=>	36598,
		1223	=>	36601,
		1224	=>	36604,
		1225	=>	36607,
		1226	=>	36610,
		1227	=>	36613,
		1228	=>	36616,
		1229	=>	36620,
		1230	=>	36623,
		1231	=>	36626,
		1232	=>	36629,
		1233	=>	36632,
		1234	=>	36635,
		1235	=>	36638,
		1236	=>	36641,
		1237	=>	36644,
		1238	=>	36648,
		1239	=>	36651,
		1240	=>	36654,
		1241	=>	36657,
		1242	=>	36660,
		1243	=>	36663,
		1244	=>	36666,
		1245	=>	36669,
		1246	=>	36673,
		1247	=>	36676,
		1248	=>	36679,
		1249	=>	36682,
		1250	=>	36685,
		1251	=>	36688,
		1252	=>	36691,
		1253	=>	36694,
		1254	=>	36698,
		1255	=>	36701,
		1256	=>	36704,
		1257	=>	36707,
		1258	=>	36710,
		1259	=>	36713,
		1260	=>	36716,
		1261	=>	36719,
		1262	=>	36722,
		1263	=>	36726,
		1264	=>	36729,
		1265	=>	36732,
		1266	=>	36735,
		1267	=>	36738,
		1268	=>	36741,
		1269	=>	36744,
		1270	=>	36747,
		1271	=>	36751,
		1272	=>	36754,
		1273	=>	36757,
		1274	=>	36760,
		1275	=>	36763,
		1276	=>	36766,
		1277	=>	36769,
		1278	=>	36772,
		1279	=>	36775,
		1280	=>	36779,
		1281	=>	36782,
		1282	=>	36785,
		1283	=>	36788,
		1284	=>	36791,
		1285	=>	36794,
		1286	=>	36797,
		1287	=>	36800,
		1288	=>	36804,
		1289	=>	36807,
		1290	=>	36810,
		1291	=>	36813,
		1292	=>	36816,
		1293	=>	36819,
		1294	=>	36822,
		1295	=>	36825,
		1296	=>	36828,
		1297	=>	36832,
		1298	=>	36835,
		1299	=>	36838,
		1300	=>	36841,
		1301	=>	36844,
		1302	=>	36847,
		1303	=>	36850,
		1304	=>	36853,
		1305	=>	36857,
		1306	=>	36860,
		1307	=>	36863,
		1308	=>	36866,
		1309	=>	36869,
		1310	=>	36872,
		1311	=>	36875,
		1312	=>	36878,
		1313	=>	36881,
		1314	=>	36885,
		1315	=>	36888,
		1316	=>	36891,
		1317	=>	36894,
		1318	=>	36897,
		1319	=>	36900,
		1320	=>	36903,
		1321	=>	36906,
		1322	=>	36910,
		1323	=>	36913,
		1324	=>	36916,
		1325	=>	36919,
		1326	=>	36922,
		1327	=>	36925,
		1328	=>	36928,
		1329	=>	36931,
		1330	=>	36934,
		1331	=>	36938,
		1332	=>	36941,
		1333	=>	36944,
		1334	=>	36947,
		1335	=>	36950,
		1336	=>	36953,
		1337	=>	36956,
		1338	=>	36959,
		1339	=>	36962,
		1340	=>	36966,
		1341	=>	36969,
		1342	=>	36972,
		1343	=>	36975,
		1344	=>	36978,
		1345	=>	36981,
		1346	=>	36984,
		1347	=>	36987,
		1348	=>	36991,
		1349	=>	36994,
		1350	=>	36997,
		1351	=>	37000,
		1352	=>	37003,
		1353	=>	37006,
		1354	=>	37009,
		1355	=>	37012,
		1356	=>	37015,
		1357	=>	37019,
		1358	=>	37022,
		1359	=>	37025,
		1360	=>	37028,
		1361	=>	37031,
		1362	=>	37034,
		1363	=>	37037,
		1364	=>	37040,
		1365	=>	37043,
		1366	=>	37047,
		1367	=>	37050,
		1368	=>	37053,
		1369	=>	37056,
		1370	=>	37059,
		1371	=>	37062,
		1372	=>	37065,
		1373	=>	37068,
		1374	=>	37072,
		1375	=>	37075,
		1376	=>	37078,
		1377	=>	37081,
		1378	=>	37084,
		1379	=>	37087,
		1380	=>	37090,
		1381	=>	37093,
		1382	=>	37096,
		1383	=>	37100,
		1384	=>	37103,
		1385	=>	37106,
		1386	=>	37109,
		1387	=>	37112,
		1388	=>	37115,
		1389	=>	37118,
		1390	=>	37121,
		1391	=>	37124,
		1392	=>	37128,
		1393	=>	37131,
		1394	=>	37134,
		1395	=>	37137,
		1396	=>	37140,
		1397	=>	37143,
		1398	=>	37146,
		1399	=>	37149,
		1400	=>	37152,
		1401	=>	37156,
		1402	=>	37159,
		1403	=>	37162,
		1404	=>	37165,
		1405	=>	37168,
		1406	=>	37171,
		1407	=>	37174,
		1408	=>	37177,
		1409	=>	37180,
		1410	=>	37184,
		1411	=>	37187,
		1412	=>	37190,
		1413	=>	37193,
		1414	=>	37196,
		1415	=>	37199,
		1416	=>	37202,
		1417	=>	37205,
		1418	=>	37209,
		1419	=>	37212,
		1420	=>	37215,
		1421	=>	37218,
		1422	=>	37221,
		1423	=>	37224,
		1424	=>	37227,
		1425	=>	37230,
		1426	=>	37233,
		1427	=>	37237,
		1428	=>	37240,
		1429	=>	37243,
		1430	=>	37246,
		1431	=>	37249,
		1432	=>	37252,
		1433	=>	37255,
		1434	=>	37258,
		1435	=>	37261,
		1436	=>	37265,
		1437	=>	37268,
		1438	=>	37271,
		1439	=>	37274,
		1440	=>	37277,
		1441	=>	37280,
		1442	=>	37283,
		1443	=>	37286,
		1444	=>	37289,
		1445	=>	37293,
		1446	=>	37296,
		1447	=>	37299,
		1448	=>	37302,
		1449	=>	37305,
		1450	=>	37308,
		1451	=>	37311,
		1452	=>	37314,
		1453	=>	37317,
		1454	=>	37321,
		1455	=>	37324,
		1456	=>	37327,
		1457	=>	37330,
		1458	=>	37333,
		1459	=>	37336,
		1460	=>	37339,
		1461	=>	37342,
		1462	=>	37345,
		1463	=>	37349,
		1464	=>	37352,
		1465	=>	37355,
		1466	=>	37358,
		1467	=>	37361,
		1468	=>	37364,
		1469	=>	37367,
		1470	=>	37370,
		1471	=>	37373,
		1472	=>	37377,
		1473	=>	37380,
		1474	=>	37383,
		1475	=>	37386,
		1476	=>	37389,
		1477	=>	37392,
		1478	=>	37395,
		1479	=>	37398,
		1480	=>	37401,
		1481	=>	37405,
		1482	=>	37408,
		1483	=>	37411,
		1484	=>	37414,
		1485	=>	37417,
		1486	=>	37420,
		1487	=>	37423,
		1488	=>	37426,
		1489	=>	37429,
		1490	=>	37432,
		1491	=>	37436,
		1492	=>	37439,
		1493	=>	37442,
		1494	=>	37445,
		1495	=>	37448,
		1496	=>	37451,
		1497	=>	37454,
		1498	=>	37457,
		1499	=>	37460,
		1500	=>	37464,
		1501	=>	37467,
		1502	=>	37470,
		1503	=>	37473,
		1504	=>	37476,
		1505	=>	37479,
		1506	=>	37482,
		1507	=>	37485,
		1508	=>	37488,
		1509	=>	37492,
		1510	=>	37495,
		1511	=>	37498,
		1512	=>	37501,
		1513	=>	37504,
		1514	=>	37507,
		1515	=>	37510,
		1516	=>	37513,
		1517	=>	37516,
		1518	=>	37520,
		1519	=>	37523,
		1520	=>	37526,
		1521	=>	37529,
		1522	=>	37532,
		1523	=>	37535,
		1524	=>	37538,
		1525	=>	37541,
		1526	=>	37544,
		1527	=>	37548,
		1528	=>	37551,
		1529	=>	37554,
		1530	=>	37557,
		1531	=>	37560,
		1532	=>	37563,
		1533	=>	37566,
		1534	=>	37569,
		1535	=>	37572,
		1536	=>	37575,
		1537	=>	37579,
		1538	=>	37582,
		1539	=>	37585,
		1540	=>	37588,
		1541	=>	37591,
		1542	=>	37594,
		1543	=>	37597,
		1544	=>	37600,
		1545	=>	37603,
		1546	=>	37607,
		1547	=>	37610,
		1548	=>	37613,
		1549	=>	37616,
		1550	=>	37619,
		1551	=>	37622,
		1552	=>	37625,
		1553	=>	37628,
		1554	=>	37631,
		1555	=>	37635,
		1556	=>	37638,
		1557	=>	37641,
		1558	=>	37644,
		1559	=>	37647,
		1560	=>	37650,
		1561	=>	37653,
		1562	=>	37656,
		1563	=>	37659,
		1564	=>	37662,
		1565	=>	37666,
		1566	=>	37669,
		1567	=>	37672,
		1568	=>	37675,
		1569	=>	37678,
		1570	=>	37681,
		1571	=>	37684,
		1572	=>	37687,
		1573	=>	37690,
		1574	=>	37694,
		1575	=>	37697,
		1576	=>	37700,
		1577	=>	37703,
		1578	=>	37706,
		1579	=>	37709,
		1580	=>	37712,
		1581	=>	37715,
		1582	=>	37718,
		1583	=>	37721,
		1584	=>	37725,
		1585	=>	37728,
		1586	=>	37731,
		1587	=>	37734,
		1588	=>	37737,
		1589	=>	37740,
		1590	=>	37743,
		1591	=>	37746,
		1592	=>	37749,
		1593	=>	37753,
		1594	=>	37756,
		1595	=>	37759,
		1596	=>	37762,
		1597	=>	37765,
		1598	=>	37768,
		1599	=>	37771,
		1600	=>	37774,
		1601	=>	37777,
		1602	=>	37780,
		1603	=>	37784,
		1604	=>	37787,
		1605	=>	37790,
		1606	=>	37793,
		1607	=>	37796,
		1608	=>	37799,
		1609	=>	37802,
		1610	=>	37805,
		1611	=>	37808,
		1612	=>	37812,
		1613	=>	37815,
		1614	=>	37818,
		1615	=>	37821,
		1616	=>	37824,
		1617	=>	37827,
		1618	=>	37830,
		1619	=>	37833,
		1620	=>	37836,
		1621	=>	37839,
		1622	=>	37843,
		1623	=>	37846,
		1624	=>	37849,
		1625	=>	37852,
		1626	=>	37855,
		1627	=>	37858,
		1628	=>	37861,
		1629	=>	37864,
		1630	=>	37867,
		1631	=>	37871,
		1632	=>	37874,
		1633	=>	37877,
		1634	=>	37880,
		1635	=>	37883,
		1636	=>	37886,
		1637	=>	37889,
		1638	=>	37892,
		1639	=>	37895,
		1640	=>	37898,
		1641	=>	37902,
		1642	=>	37905,
		1643	=>	37908,
		1644	=>	37911,
		1645	=>	37914,
		1646	=>	37917,
		1647	=>	37920,
		1648	=>	37923,
		1649	=>	37926,
		1650	=>	37929,
		1651	=>	37933,
		1652	=>	37936,
		1653	=>	37939,
		1654	=>	37942,
		1655	=>	37945,
		1656	=>	37948,
		1657	=>	37951,
		1658	=>	37954,
		1659	=>	37957,
		1660	=>	37960,
		1661	=>	37964,
		1662	=>	37967,
		1663	=>	37970,
		1664	=>	37973,
		1665	=>	37976,
		1666	=>	37979,
		1667	=>	37982,
		1668	=>	37985,
		1669	=>	37988,
		1670	=>	37991,
		1671	=>	37995,
		1672	=>	37998,
		1673	=>	38001,
		1674	=>	38004,
		1675	=>	38007,
		1676	=>	38010,
		1677	=>	38013,
		1678	=>	38016,
		1679	=>	38019,
		1680	=>	38023,
		1681	=>	38026,
		1682	=>	38029,
		1683	=>	38032,
		1684	=>	38035,
		1685	=>	38038,
		1686	=>	38041,
		1687	=>	38044,
		1688	=>	38047,
		1689	=>	38050,
		1690	=>	38054,
		1691	=>	38057,
		1692	=>	38060,
		1693	=>	38063,
		1694	=>	38066,
		1695	=>	38069,
		1696	=>	38072,
		1697	=>	38075,
		1698	=>	38078,
		1699	=>	38081,
		1700	=>	38085,
		1701	=>	38088,
		1702	=>	38091,
		1703	=>	38094,
		1704	=>	38097,
		1705	=>	38100,
		1706	=>	38103,
		1707	=>	38106,
		1708	=>	38109,
		1709	=>	38112,
		1710	=>	38116,
		1711	=>	38119,
		1712	=>	38122,
		1713	=>	38125,
		1714	=>	38128,
		1715	=>	38131,
		1716	=>	38134,
		1717	=>	38137,
		1718	=>	38140,
		1719	=>	38143,
		1720	=>	38147,
		1721	=>	38150,
		1722	=>	38153,
		1723	=>	38156,
		1724	=>	38159,
		1725	=>	38162,
		1726	=>	38165,
		1727	=>	38168,
		1728	=>	38171,
		1729	=>	38174,
		1730	=>	38177,
		1731	=>	38181,
		1732	=>	38184,
		1733	=>	38187,
		1734	=>	38190,
		1735	=>	38193,
		1736	=>	38196,
		1737	=>	38199,
		1738	=>	38202,
		1739	=>	38205,
		1740	=>	38208,
		1741	=>	38212,
		1742	=>	38215,
		1743	=>	38218,
		1744	=>	38221,
		1745	=>	38224,
		1746	=>	38227,
		1747	=>	38230,
		1748	=>	38233,
		1749	=>	38236,
		1750	=>	38239,
		1751	=>	38243,
		1752	=>	38246,
		1753	=>	38249,
		1754	=>	38252,
		1755	=>	38255,
		1756	=>	38258,
		1757	=>	38261,
		1758	=>	38264,
		1759	=>	38267,
		1760	=>	38270,
		1761	=>	38274,
		1762	=>	38277,
		1763	=>	38280,
		1764	=>	38283,
		1765	=>	38286,
		1766	=>	38289,
		1767	=>	38292,
		1768	=>	38295,
		1769	=>	38298,
		1770	=>	38301,
		1771	=>	38304,
		1772	=>	38308,
		1773	=>	38311,
		1774	=>	38314,
		1775	=>	38317,
		1776	=>	38320,
		1777	=>	38323,
		1778	=>	38326,
		1779	=>	38329,
		1780	=>	38332,
		1781	=>	38335,
		1782	=>	38339,
		1783	=>	38342,
		1784	=>	38345,
		1785	=>	38348,
		1786	=>	38351,
		1787	=>	38354,
		1788	=>	38357,
		1789	=>	38360,
		1790	=>	38363,
		1791	=>	38366,
		1792	=>	38369,
		1793	=>	38373,
		1794	=>	38376,
		1795	=>	38379,
		1796	=>	38382,
		1797	=>	38385,
		1798	=>	38388,
		1799	=>	38391,
		1800	=>	38394,
		1801	=>	38397,
		1802	=>	38400,
		1803	=>	38404,
		1804	=>	38407,
		1805	=>	38410,
		1806	=>	38413,
		1807	=>	38416,
		1808	=>	38419,
		1809	=>	38422,
		1810	=>	38425,
		1811	=>	38428,
		1812	=>	38431,
		1813	=>	38434,
		1814	=>	38438,
		1815	=>	38441,
		1816	=>	38444,
		1817	=>	38447,
		1818	=>	38450,
		1819	=>	38453,
		1820	=>	38456,
		1821	=>	38459,
		1822	=>	38462,
		1823	=>	38465,
		1824	=>	38469,
		1825	=>	38472,
		1826	=>	38475,
		1827	=>	38478,
		1828	=>	38481,
		1829	=>	38484,
		1830	=>	38487,
		1831	=>	38490,
		1832	=>	38493,
		1833	=>	38496,
		1834	=>	38499,
		1835	=>	38503,
		1836	=>	38506,
		1837	=>	38509,
		1838	=>	38512,
		1839	=>	38515,
		1840	=>	38518,
		1841	=>	38521,
		1842	=>	38524,
		1843	=>	38527,
		1844	=>	38530,
		1845	=>	38533,
		1846	=>	38537,
		1847	=>	38540,
		1848	=>	38543,
		1849	=>	38546,
		1850	=>	38549,
		1851	=>	38552,
		1852	=>	38555,
		1853	=>	38558,
		1854	=>	38561,
		1855	=>	38564,
		1856	=>	38567,
		1857	=>	38571,
		1858	=>	38574,
		1859	=>	38577,
		1860	=>	38580,
		1861	=>	38583,
		1862	=>	38586,
		1863	=>	38589,
		1864	=>	38592,
		1865	=>	38595,
		1866	=>	38598,
		1867	=>	38601,
		1868	=>	38605,
		1869	=>	38608,
		1870	=>	38611,
		1871	=>	38614,
		1872	=>	38617,
		1873	=>	38620,
		1874	=>	38623,
		1875	=>	38626,
		1876	=>	38629,
		1877	=>	38632,
		1878	=>	38635,
		1879	=>	38639,
		1880	=>	38642,
		1881	=>	38645,
		1882	=>	38648,
		1883	=>	38651,
		1884	=>	38654,
		1885	=>	38657,
		1886	=>	38660,
		1887	=>	38663,
		1888	=>	38666,
		1889	=>	38669,
		1890	=>	38673,
		1891	=>	38676,
		1892	=>	38679,
		1893	=>	38682,
		1894	=>	38685,
		1895	=>	38688,
		1896	=>	38691,
		1897	=>	38694,
		1898	=>	38697,
		1899	=>	38700,
		1900	=>	38703,
		1901	=>	38707,
		1902	=>	38710,
		1903	=>	38713,
		1904	=>	38716,
		1905	=>	38719,
		1906	=>	38722,
		1907	=>	38725,
		1908	=>	38728,
		1909	=>	38731,
		1910	=>	38734,
		1911	=>	38737,
		1912	=>	38741,
		1913	=>	38744,
		1914	=>	38747,
		1915	=>	38750,
		1916	=>	38753,
		1917	=>	38756,
		1918	=>	38759,
		1919	=>	38762,
		1920	=>	38765,
		1921	=>	38768,
		1922	=>	38771,
		1923	=>	38775,
		1924	=>	38778,
		1925	=>	38781,
		1926	=>	38784,
		1927	=>	38787,
		1928	=>	38790,
		1929	=>	38793,
		1930	=>	38796,
		1931	=>	38799,
		1932	=>	38802,
		1933	=>	38805,
		1934	=>	38808,
		1935	=>	38812,
		1936	=>	38815,
		1937	=>	38818,
		1938	=>	38821,
		1939	=>	38824,
		1940	=>	38827,
		1941	=>	38830,
		1942	=>	38833,
		1943	=>	38836,
		1944	=>	38839,
		1945	=>	38842,
		1946	=>	38846,
		1947	=>	38849,
		1948	=>	38852,
		1949	=>	38855,
		1950	=>	38858,
		1951	=>	38861,
		1952	=>	38864,
		1953	=>	38867,
		1954	=>	38870,
		1955	=>	38873,
		1956	=>	38876,
		1957	=>	38879,
		1958	=>	38883,
		1959	=>	38886,
		1960	=>	38889,
		1961	=>	38892,
		1962	=>	38895,
		1963	=>	38898,
		1964	=>	38901,
		1965	=>	38904,
		1966	=>	38907,
		1967	=>	38910,
		1968	=>	38913,
		1969	=>	38917,
		1970	=>	38920,
		1971	=>	38923,
		1972	=>	38926,
		1973	=>	38929,
		1974	=>	38932,
		1975	=>	38935,
		1976	=>	38938,
		1977	=>	38941,
		1978	=>	38944,
		1979	=>	38947,
		1980	=>	38950,
		1981	=>	38954,
		1982	=>	38957,
		1983	=>	38960,
		1984	=>	38963,
		1985	=>	38966,
		1986	=>	38969,
		1987	=>	38972,
		1988	=>	38975,
		1989	=>	38978,
		1990	=>	38981,
		1991	=>	38984,
		1992	=>	38987,
		1993	=>	38991,
		1994	=>	38994,
		1995	=>	38997,
		1996	=>	39000,
		1997	=>	39003,
		1998	=>	39006,
		1999	=>	39009,
		2000	=>	39012,
		2001	=>	39015,
		2002	=>	39018,
		2003	=>	39021,
		2004	=>	39024,
		2005	=>	39028,
		2006	=>	39031,
		2007	=>	39034,
		2008	=>	39037,
		2009	=>	39040,
		2010	=>	39043,
		2011	=>	39046,
		2012	=>	39049,
		2013	=>	39052,
		2014	=>	39055,
		2015	=>	39058,
		2016	=>	39061,
		2017	=>	39065,
		2018	=>	39068,
		2019	=>	39071,
		2020	=>	39074,
		2021	=>	39077,
		2022	=>	39080,
		2023	=>	39083,
		2024	=>	39086,
		2025	=>	39089,
		2026	=>	39092,
		2027	=>	39095,
		2028	=>	39098,
		2029	=>	39102,
		2030	=>	39105,
		2031	=>	39108,
		2032	=>	39111,
		2033	=>	39114,
		2034	=>	39117,
		2035	=>	39120,
		2036	=>	39123,
		2037	=>	39126,
		2038	=>	39129,
		2039	=>	39132,
		2040	=>	39135,
		2041	=>	39139,
		2042	=>	39142,
		2043	=>	39145,
		2044	=>	39148,
		2045	=>	39151,
		2046	=>	39154,
		2047	=>	39157,
		2048	=>	39160,
		2049	=>	39163,
		2050	=>	39166,
		2051	=>	39169,
		2052	=>	39172,
		2053	=>	39176,
		2054	=>	39179,
		2055	=>	39182,
		2056	=>	39185,
		2057	=>	39188,
		2058	=>	39191,
		2059	=>	39194,
		2060	=>	39197,
		2061	=>	39200,
		2062	=>	39203,
		2063	=>	39206,
		2064	=>	39209,
		2065	=>	39212,
		2066	=>	39216,
		2067	=>	39219,
		2068	=>	39222,
		2069	=>	39225,
		2070	=>	39228,
		2071	=>	39231,
		2072	=>	39234,
		2073	=>	39237,
		2074	=>	39240,
		2075	=>	39243,
		2076	=>	39246,
		2077	=>	39249,
		2078	=>	39253,
		2079	=>	39256,
		2080	=>	39259,
		2081	=>	39262,
		2082	=>	39265,
		2083	=>	39268,
		2084	=>	39271,
		2085	=>	39274,
		2086	=>	39277,
		2087	=>	39280,
		2088	=>	39283,
		2089	=>	39286,
		2090	=>	39289,
		2091	=>	39293,
		2092	=>	39296,
		2093	=>	39299,
		2094	=>	39302,
		2095	=>	39305,
		2096	=>	39308,
		2097	=>	39311,
		2098	=>	39314,
		2099	=>	39317,
		2100	=>	39320,
		2101	=>	39323,
		2102	=>	39326,
		2103	=>	39329,
		2104	=>	39333,
		2105	=>	39336,
		2106	=>	39339,
		2107	=>	39342,
		2108	=>	39345,
		2109	=>	39348,
		2110	=>	39351,
		2111	=>	39354,
		2112	=>	39357,
		2113	=>	39360,
		2114	=>	39363,
		2115	=>	39366,
		2116	=>	39370,
		2117	=>	39373,
		2118	=>	39376,
		2119	=>	39379,
		2120	=>	39382,
		2121	=>	39385,
		2122	=>	39388,
		2123	=>	39391,
		2124	=>	39394,
		2125	=>	39397,
		2126	=>	39400,
		2127	=>	39403,
		2128	=>	39406,
		2129	=>	39410,
		2130	=>	39413,
		2131	=>	39416,
		2132	=>	39419,
		2133	=>	39422,
		2134	=>	39425,
		2135	=>	39428,
		2136	=>	39431,
		2137	=>	39434,
		2138	=>	39437,
		2139	=>	39440,
		2140	=>	39443,
		2141	=>	39446,
		2142	=>	39449,
		2143	=>	39453,
		2144	=>	39456,
		2145	=>	39459,
		2146	=>	39462,
		2147	=>	39465,
		2148	=>	39468,
		2149	=>	39471,
		2150	=>	39474,
		2151	=>	39477,
		2152	=>	39480,
		2153	=>	39483,
		2154	=>	39486,
		2155	=>	39489,
		2156	=>	39493,
		2157	=>	39496,
		2158	=>	39499,
		2159	=>	39502,
		2160	=>	39505,
		2161	=>	39508,
		2162	=>	39511,
		2163	=>	39514,
		2164	=>	39517,
		2165	=>	39520,
		2166	=>	39523,
		2167	=>	39526,
		2168	=>	39529,
		2169	=>	39533,
		2170	=>	39536,
		2171	=>	39539,
		2172	=>	39542,
		2173	=>	39545,
		2174	=>	39548,
		2175	=>	39551,
		2176	=>	39554,
		2177	=>	39557,
		2178	=>	39560,
		2179	=>	39563,
		2180	=>	39566,
		2181	=>	39569,
		2182	=>	39572,
		2183	=>	39576,
		2184	=>	39579,
		2185	=>	39582,
		2186	=>	39585,
		2187	=>	39588,
		2188	=>	39591,
		2189	=>	39594,
		2190	=>	39597,
		2191	=>	39600,
		2192	=>	39603,
		2193	=>	39606,
		2194	=>	39609,
		2195	=>	39612,
		2196	=>	39615,
		2197	=>	39619,
		2198	=>	39622,
		2199	=>	39625,
		2200	=>	39628,
		2201	=>	39631,
		2202	=>	39634,
		2203	=>	39637,
		2204	=>	39640,
		2205	=>	39643,
		2206	=>	39646,
		2207	=>	39649,
		2208	=>	39652,
		2209	=>	39655,
		2210	=>	39658,
		2211	=>	39662,
		2212	=>	39665,
		2213	=>	39668,
		2214	=>	39671,
		2215	=>	39674,
		2216	=>	39677,
		2217	=>	39680,
		2218	=>	39683,
		2219	=>	39686,
		2220	=>	39689,
		2221	=>	39692,
		2222	=>	39695,
		2223	=>	39698,
		2224	=>	39701,
		2225	=>	39705,
		2226	=>	39708,
		2227	=>	39711,
		2228	=>	39714,
		2229	=>	39717,
		2230	=>	39720,
		2231	=>	39723,
		2232	=>	39726,
		2233	=>	39729,
		2234	=>	39732,
		2235	=>	39735,
		2236	=>	39738,
		2237	=>	39741,
		2238	=>	39744,
		2239	=>	39748,
		2240	=>	39751,
		2241	=>	39754,
		2242	=>	39757,
		2243	=>	39760,
		2244	=>	39763,
		2245	=>	39766,
		2246	=>	39769,
		2247	=>	39772,
		2248	=>	39775,
		2249	=>	39778,
		2250	=>	39781,
		2251	=>	39784,
		2252	=>	39787,
		2253	=>	39790,
		2254	=>	39794,
		2255	=>	39797,
		2256	=>	39800,
		2257	=>	39803,
		2258	=>	39806,
		2259	=>	39809,
		2260	=>	39812,
		2261	=>	39815,
		2262	=>	39818,
		2263	=>	39821,
		2264	=>	39824,
		2265	=>	39827,
		2266	=>	39830,
		2267	=>	39833,
		2268	=>	39837,
		2269	=>	39840,
		2270	=>	39843,
		2271	=>	39846,
		2272	=>	39849,
		2273	=>	39852,
		2274	=>	39855,
		2275	=>	39858,
		2276	=>	39861,
		2277	=>	39864,
		2278	=>	39867,
		2279	=>	39870,
		2280	=>	39873,
		2281	=>	39876,
		2282	=>	39879,
		2283	=>	39883,
		2284	=>	39886,
		2285	=>	39889,
		2286	=>	39892,
		2287	=>	39895,
		2288	=>	39898,
		2289	=>	39901,
		2290	=>	39904,
		2291	=>	39907,
		2292	=>	39910,
		2293	=>	39913,
		2294	=>	39916,
		2295	=>	39919,
		2296	=>	39922,
		2297	=>	39925,
		2298	=>	39929,
		2299	=>	39932,
		2300	=>	39935,
		2301	=>	39938,
		2302	=>	39941,
		2303	=>	39944,
		2304	=>	39947,
		2305	=>	39950,
		2306	=>	39953,
		2307	=>	39956,
		2308	=>	39959,
		2309	=>	39962,
		2310	=>	39965,
		2311	=>	39968,
		2312	=>	39971,
		2313	=>	39974,
		2314	=>	39978,
		2315	=>	39981,
		2316	=>	39984,
		2317	=>	39987,
		2318	=>	39990,
		2319	=>	39993,
		2320	=>	39996,
		2321	=>	39999,
		2322	=>	40002,
		2323	=>	40005,
		2324	=>	40008,
		2325	=>	40011,
		2326	=>	40014,
		2327	=>	40017,
		2328	=>	40020,
		2329	=>	40024,
		2330	=>	40027,
		2331	=>	40030,
		2332	=>	40033,
		2333	=>	40036,
		2334	=>	40039,
		2335	=>	40042,
		2336	=>	40045,
		2337	=>	40048,
		2338	=>	40051,
		2339	=>	40054,
		2340	=>	40057,
		2341	=>	40060,
		2342	=>	40063,
		2343	=>	40066,
		2344	=>	40069,
		2345	=>	40073,
		2346	=>	40076,
		2347	=>	40079,
		2348	=>	40082,
		2349	=>	40085,
		2350	=>	40088,
		2351	=>	40091,
		2352	=>	40094,
		2353	=>	40097,
		2354	=>	40100,
		2355	=>	40103,
		2356	=>	40106,
		2357	=>	40109,
		2358	=>	40112,
		2359	=>	40115,
		2360	=>	40118,
		2361	=>	40122,
		2362	=>	40125,
		2363	=>	40128,
		2364	=>	40131,
		2365	=>	40134,
		2366	=>	40137,
		2367	=>	40140,
		2368	=>	40143,
		2369	=>	40146,
		2370	=>	40149,
		2371	=>	40152,
		2372	=>	40155,
		2373	=>	40158,
		2374	=>	40161,
		2375	=>	40164,
		2376	=>	40167,
		2377	=>	40170,
		2378	=>	40174,
		2379	=>	40177,
		2380	=>	40180,
		2381	=>	40183,
		2382	=>	40186,
		2383	=>	40189,
		2384	=>	40192,
		2385	=>	40195,
		2386	=>	40198,
		2387	=>	40201,
		2388	=>	40204,
		2389	=>	40207,
		2390	=>	40210,
		2391	=>	40213,
		2392	=>	40216,
		2393	=>	40219,
		2394	=>	40222,
		2395	=>	40226,
		2396	=>	40229,
		2397	=>	40232,
		2398	=>	40235,
		2399	=>	40238,
		2400	=>	40241,
		2401	=>	40244,
		2402	=>	40247,
		2403	=>	40250,
		2404	=>	40253,
		2405	=>	40256,
		2406	=>	40259,
		2407	=>	40262,
		2408	=>	40265,
		2409	=>	40268,
		2410	=>	40271,
		2411	=>	40274,
		2412	=>	40278,
		2413	=>	40281,
		2414	=>	40284,
		2415	=>	40287,
		2416	=>	40290,
		2417	=>	40293,
		2418	=>	40296,
		2419	=>	40299,
		2420	=>	40302,
		2421	=>	40305,
		2422	=>	40308,
		2423	=>	40311,
		2424	=>	40314,
		2425	=>	40317,
		2426	=>	40320,
		2427	=>	40323,
		2428	=>	40326,
		2429	=>	40330,
		2430	=>	40333,
		2431	=>	40336,
		2432	=>	40339,
		2433	=>	40342,
		2434	=>	40345,
		2435	=>	40348,
		2436	=>	40351,
		2437	=>	40354,
		2438	=>	40357,
		2439	=>	40360,
		2440	=>	40363,
		2441	=>	40366,
		2442	=>	40369,
		2443	=>	40372,
		2444	=>	40375,
		2445	=>	40378,
		2446	=>	40381,
		2447	=>	40385,
		2448	=>	40388,
		2449	=>	40391,
		2450	=>	40394,
		2451	=>	40397,
		2452	=>	40400,
		2453	=>	40403,
		2454	=>	40406,
		2455	=>	40409,
		2456	=>	40412,
		2457	=>	40415,
		2458	=>	40418,
		2459	=>	40421,
		2460	=>	40424,
		2461	=>	40427,
		2462	=>	40430,
		2463	=>	40433,
		2464	=>	40436,
		2465	=>	40440,
		2466	=>	40443,
		2467	=>	40446,
		2468	=>	40449,
		2469	=>	40452,
		2470	=>	40455,
		2471	=>	40458,
		2472	=>	40461,
		2473	=>	40464,
		2474	=>	40467,
		2475	=>	40470,
		2476	=>	40473,
		2477	=>	40476,
		2478	=>	40479,
		2479	=>	40482,
		2480	=>	40485,
		2481	=>	40488,
		2482	=>	40491,
		2483	=>	40494,
		2484	=>	40498,
		2485	=>	40501,
		2486	=>	40504,
		2487	=>	40507,
		2488	=>	40510,
		2489	=>	40513,
		2490	=>	40516,
		2491	=>	40519,
		2492	=>	40522,
		2493	=>	40525,
		2494	=>	40528,
		2495	=>	40531,
		2496	=>	40534,
		2497	=>	40537,
		2498	=>	40540,
		2499	=>	40543,
		2500	=>	40546,
		2501	=>	40549,
		2502	=>	40552,
		2503	=>	40556,
		2504	=>	40559,
		2505	=>	40562,
		2506	=>	40565,
		2507	=>	40568,
		2508	=>	40571,
		2509	=>	40574,
		2510	=>	40577,
		2511	=>	40580,
		2512	=>	40583,
		2513	=>	40586,
		2514	=>	40589,
		2515	=>	40592,
		2516	=>	40595,
		2517	=>	40598,
		2518	=>	40601,
		2519	=>	40604,
		2520	=>	40607,
		2521	=>	40610,
		2522	=>	40613,
		2523	=>	40617,
		2524	=>	40620,
		2525	=>	40623,
		2526	=>	40626,
		2527	=>	40629,
		2528	=>	40632,
		2529	=>	40635,
		2530	=>	40638,
		2531	=>	40641,
		2532	=>	40644,
		2533	=>	40647,
		2534	=>	40650,
		2535	=>	40653,
		2536	=>	40656,
		2537	=>	40659,
		2538	=>	40662,
		2539	=>	40665,
		2540	=>	40668,
		2541	=>	40671,
		2542	=>	40674,
		2543	=>	40678,
		2544	=>	40681,
		2545	=>	40684,
		2546	=>	40687,
		2547	=>	40690,
		2548	=>	40693,
		2549	=>	40696,
		2550	=>	40699,
		2551	=>	40702,
		2552	=>	40705,
		2553	=>	40708,
		2554	=>	40711,
		2555	=>	40714,
		2556	=>	40717,
		2557	=>	40720,
		2558	=>	40723,
		2559	=>	40726,
		2560	=>	40729,
		2561	=>	40732,
		2562	=>	40735,
		2563	=>	40738,
		2564	=>	40742,
		2565	=>	40745,
		2566	=>	40748,
		2567	=>	40751,
		2568	=>	40754,
		2569	=>	40757,
		2570	=>	40760,
		2571	=>	40763,
		2572	=>	40766,
		2573	=>	40769,
		2574	=>	40772,
		2575	=>	40775,
		2576	=>	40778,
		2577	=>	40781,
		2578	=>	40784,
		2579	=>	40787,
		2580	=>	40790,
		2581	=>	40793,
		2582	=>	40796,
		2583	=>	40799,
		2584	=>	40802,
		2585	=>	40806,
		2586	=>	40809,
		2587	=>	40812,
		2588	=>	40815,
		2589	=>	40818,
		2590	=>	40821,
		2591	=>	40824,
		2592	=>	40827,
		2593	=>	40830,
		2594	=>	40833,
		2595	=>	40836,
		2596	=>	40839,
		2597	=>	40842,
		2598	=>	40845,
		2599	=>	40848,
		2600	=>	40851,
		2601	=>	40854,
		2602	=>	40857,
		2603	=>	40860,
		2604	=>	40863,
		2605	=>	40866,
		2606	=>	40869,
		2607	=>	40872,
		2608	=>	40876,
		2609	=>	40879,
		2610	=>	40882,
		2611	=>	40885,
		2612	=>	40888,
		2613	=>	40891,
		2614	=>	40894,
		2615	=>	40897,
		2616	=>	40900,
		2617	=>	40903,
		2618	=>	40906,
		2619	=>	40909,
		2620	=>	40912,
		2621	=>	40915,
		2622	=>	40918,
		2623	=>	40921,
		2624	=>	40924,
		2625	=>	40927,
		2626	=>	40930,
		2627	=>	40933,
		2628	=>	40936,
		2629	=>	40939,
		2630	=>	40942,
		2631	=>	40946,
		2632	=>	40949,
		2633	=>	40952,
		2634	=>	40955,
		2635	=>	40958,
		2636	=>	40961,
		2637	=>	40964,
		2638	=>	40967,
		2639	=>	40970,
		2640	=>	40973,
		2641	=>	40976,
		2642	=>	40979,
		2643	=>	40982,
		2644	=>	40985,
		2645	=>	40988,
		2646	=>	40991,
		2647	=>	40994,
		2648	=>	40997,
		2649	=>	41000,
		2650	=>	41003,
		2651	=>	41006,
		2652	=>	41009,
		2653	=>	41012,
		2654	=>	41015,
		2655	=>	41019,
		2656	=>	41022,
		2657	=>	41025,
		2658	=>	41028,
		2659	=>	41031,
		2660	=>	41034,
		2661	=>	41037,
		2662	=>	41040,
		2663	=>	41043,
		2664	=>	41046,
		2665	=>	41049,
		2666	=>	41052,
		2667	=>	41055,
		2668	=>	41058,
		2669	=>	41061,
		2670	=>	41064,
		2671	=>	41067,
		2672	=>	41070,
		2673	=>	41073,
		2674	=>	41076,
		2675	=>	41079,
		2676	=>	41082,
		2677	=>	41085,
		2678	=>	41088,
		2679	=>	41091,
		2680	=>	41095,
		2681	=>	41098,
		2682	=>	41101,
		2683	=>	41104,
		2684	=>	41107,
		2685	=>	41110,
		2686	=>	41113,
		2687	=>	41116,
		2688	=>	41119,
		2689	=>	41122,
		2690	=>	41125,
		2691	=>	41128,
		2692	=>	41131,
		2693	=>	41134,
		2694	=>	41137,
		2695	=>	41140,
		2696	=>	41143,
		2697	=>	41146,
		2698	=>	41149,
		2699	=>	41152,
		2700	=>	41155,
		2701	=>	41158,
		2702	=>	41161,
		2703	=>	41164,
		2704	=>	41167,
		2705	=>	41170,
		2706	=>	41173,
		2707	=>	41177,
		2708	=>	41180,
		2709	=>	41183,
		2710	=>	41186,
		2711	=>	41189,
		2712	=>	41192,
		2713	=>	41195,
		2714	=>	41198,
		2715	=>	41201,
		2716	=>	41204,
		2717	=>	41207,
		2718	=>	41210,
		2719	=>	41213,
		2720	=>	41216,
		2721	=>	41219,
		2722	=>	41222,
		2723	=>	41225,
		2724	=>	41228,
		2725	=>	41231,
		2726	=>	41234,
		2727	=>	41237,
		2728	=>	41240,
		2729	=>	41243,
		2730	=>	41246,
		2731	=>	41249,
		2732	=>	41252,
		2733	=>	41255,
		2734	=>	41258,
		2735	=>	41262,
		2736	=>	41265,
		2737	=>	41268,
		2738	=>	41271,
		2739	=>	41274,
		2740	=>	41277,
		2741	=>	41280,
		2742	=>	41283,
		2743	=>	41286,
		2744	=>	41289,
		2745	=>	41292,
		2746	=>	41295,
		2747	=>	41298,
		2748	=>	41301,
		2749	=>	41304,
		2750	=>	41307,
		2751	=>	41310,
		2752	=>	41313,
		2753	=>	41316,
		2754	=>	41319,
		2755	=>	41322,
		2756	=>	41325,
		2757	=>	41328,
		2758	=>	41331,
		2759	=>	41334,
		2760	=>	41337,
		2761	=>	41340,
		2762	=>	41343,
		2763	=>	41346,
		2764	=>	41349,
		2765	=>	41352,
		2766	=>	41356,
		2767	=>	41359,
		2768	=>	41362,
		2769	=>	41365,
		2770	=>	41368,
		2771	=>	41371,
		2772	=>	41374,
		2773	=>	41377,
		2774	=>	41380,
		2775	=>	41383,
		2776	=>	41386,
		2777	=>	41389,
		2778	=>	41392,
		2779	=>	41395,
		2780	=>	41398,
		2781	=>	41401,
		2782	=>	41404,
		2783	=>	41407,
		2784	=>	41410,
		2785	=>	41413,
		2786	=>	41416,
		2787	=>	41419,
		2788	=>	41422,
		2789	=>	41425,
		2790	=>	41428,
		2791	=>	41431,
		2792	=>	41434,
		2793	=>	41437,
		2794	=>	41440,
		2795	=>	41443,
		2796	=>	41446,
		2797	=>	41449,
		2798	=>	41452,
		2799	=>	41456,
		2800	=>	41459,
		2801	=>	41462,
		2802	=>	41465,
		2803	=>	41468,
		2804	=>	41471,
		2805	=>	41474,
		2806	=>	41477,
		2807	=>	41480,
		2808	=>	41483,
		2809	=>	41486,
		2810	=>	41489,
		2811	=>	41492,
		2812	=>	41495,
		2813	=>	41498,
		2814	=>	41501,
		2815	=>	41504,
		2816	=>	41507,
		2817	=>	41510,
		2818	=>	41513,
		2819	=>	41516,
		2820	=>	41519,
		2821	=>	41522,
		2822	=>	41525,
		2823	=>	41528,
		2824	=>	41531,
		2825	=>	41534,
		2826	=>	41537,
		2827	=>	41540,
		2828	=>	41543,
		2829	=>	41546,
		2830	=>	41549,
		2831	=>	41552,
		2832	=>	41555,
		2833	=>	41558,
		2834	=>	41561,
		2835	=>	41565,
		2836	=>	41568,
		2837	=>	41571,
		2838	=>	41574,
		2839	=>	41577,
		2840	=>	41580,
		2841	=>	41583,
		2842	=>	41586,
		2843	=>	41589,
		2844	=>	41592,
		2845	=>	41595,
		2846	=>	41598,
		2847	=>	41601,
		2848	=>	41604,
		2849	=>	41607,
		2850	=>	41610,
		2851	=>	41613,
		2852	=>	41616,
		2853	=>	41619,
		2854	=>	41622,
		2855	=>	41625,
		2856	=>	41628,
		2857	=>	41631,
		2858	=>	41634,
		2859	=>	41637,
		2860	=>	41640,
		2861	=>	41643,
		2862	=>	41646,
		2863	=>	41649,
		2864	=>	41652,
		2865	=>	41655,
		2866	=>	41658,
		2867	=>	41661,
		2868	=>	41664,
		2869	=>	41667,
		2870	=>	41670,
		2871	=>	41673,
		2872	=>	41676,
		2873	=>	41679,
		2874	=>	41682,
		2875	=>	41686,
		2876	=>	41689,
		2877	=>	41692,
		2878	=>	41695,
		2879	=>	41698,
		2880	=>	41701,
		2881	=>	41704,
		2882	=>	41707,
		2883	=>	41710,
		2884	=>	41713,
		2885	=>	41716,
		2886	=>	41719,
		2887	=>	41722,
		2888	=>	41725,
		2889	=>	41728,
		2890	=>	41731,
		2891	=>	41734,
		2892	=>	41737,
		2893	=>	41740,
		2894	=>	41743,
		2895	=>	41746,
		2896	=>	41749,
		2897	=>	41752,
		2898	=>	41755,
		2899	=>	41758,
		2900	=>	41761,
		2901	=>	41764,
		2902	=>	41767,
		2903	=>	41770,
		2904	=>	41773,
		2905	=>	41776,
		2906	=>	41779,
		2907	=>	41782,
		2908	=>	41785,
		2909	=>	41788,
		2910	=>	41791,
		2911	=>	41794,
		2912	=>	41797,
		2913	=>	41800,
		2914	=>	41803,
		2915	=>	41806,
		2916	=>	41809,
		2917	=>	41812,
		2918	=>	41815,
		2919	=>	41818,
		2920	=>	41821,
		2921	=>	41824,
		2922	=>	41827,
		2923	=>	41831,
		2924	=>	41834,
		2925	=>	41837,
		2926	=>	41840,
		2927	=>	41843,
		2928	=>	41846,
		2929	=>	41849,
		2930	=>	41852,
		2931	=>	41855,
		2932	=>	41858,
		2933	=>	41861,
		2934	=>	41864,
		2935	=>	41867,
		2936	=>	41870,
		2937	=>	41873,
		2938	=>	41876,
		2939	=>	41879,
		2940	=>	41882,
		2941	=>	41885,
		2942	=>	41888,
		2943	=>	41891,
		2944	=>	41894,
		2945	=>	41897,
		2946	=>	41900,
		2947	=>	41903,
		2948	=>	41906,
		2949	=>	41909,
		2950	=>	41912,
		2951	=>	41915,
		2952	=>	41918,
		2953	=>	41921,
		2954	=>	41924,
		2955	=>	41927,
		2956	=>	41930,
		2957	=>	41933,
		2958	=>	41936,
		2959	=>	41939,
		2960	=>	41942,
		2961	=>	41945,
		2962	=>	41948,
		2963	=>	41951,
		2964	=>	41954,
		2965	=>	41957,
		2966	=>	41960,
		2967	=>	41963,
		2968	=>	41966,
		2969	=>	41969,
		2970	=>	41972,
		2971	=>	41975,
		2972	=>	41978,
		2973	=>	41981,
		2974	=>	41984,
		2975	=>	41987,
		2976	=>	41990,
		2977	=>	41993,
		2978	=>	41996,
		2979	=>	41999,
		2980	=>	42002,
		2981	=>	42005,
		2982	=>	42008,
		2983	=>	42012,
		2984	=>	42015,
		2985	=>	42018,
		2986	=>	42021,
		2987	=>	42024,
		2988	=>	42027,
		2989	=>	42030,
		2990	=>	42033,
		2991	=>	42036,
		2992	=>	42039,
		2993	=>	42042,
		2994	=>	42045,
		2995	=>	42048,
		2996	=>	42051,
		2997	=>	42054,
		2998	=>	42057,
		2999	=>	42060,
		3000	=>	42063,
		3001	=>	42066,
		3002	=>	42069,
		3003	=>	42072,
		3004	=>	42075,
		3005	=>	42078,
		3006	=>	42081,
		3007	=>	42084,
		3008	=>	42087,
		3009	=>	42090,
		3010	=>	42093,
		3011	=>	42096,
		3012	=>	42099,
		3013	=>	42102,
		3014	=>	42105,
		3015	=>	42108,
		3016	=>	42111,
		3017	=>	42114,
		3018	=>	42117,
		3019	=>	42120,
		3020	=>	42123,
		3021	=>	42126,
		3022	=>	42129,
		3023	=>	42132,
		3024	=>	42135,
		3025	=>	42138,
		3026	=>	42141,
		3027	=>	42144,
		3028	=>	42147,
		3029	=>	42150,
		3030	=>	42153,
		3031	=>	42156,
		3032	=>	42159,
		3033	=>	42162,
		3034	=>	42165,
		3035	=>	42168,
		3036	=>	42171,
		3037	=>	42174,
		3038	=>	42177,
		3039	=>	42180,
		3040	=>	42183,
		3041	=>	42186,
		3042	=>	42189,
		3043	=>	42192,
		3044	=>	42195,
		3045	=>	42198,
		3046	=>	42201,
		3047	=>	42204,
		3048	=>	42207,
		3049	=>	42210,
		3050	=>	42213,
		3051	=>	42216,
		3052	=>	42219,
		3053	=>	42222,
		3054	=>	42225,
		3055	=>	42228,
		3056	=>	42231,
		3057	=>	42234,
		3058	=>	42237,
		3059	=>	42240,
		3060	=>	42243,
		3061	=>	42246,
		3062	=>	42249,
		3063	=>	42252,
		3064	=>	42255,
		3065	=>	42258,
		3066	=>	42261,
		3067	=>	42264,
		3068	=>	42267,
		3069	=>	42270,
		3070	=>	42273,
		3071	=>	42276,
		3072	=>	42279,
		3073	=>	42282,
		3074	=>	42285,
		3075	=>	42288,
		3076	=>	42291,
		3077	=>	42294,
		3078	=>	42297,
		3079	=>	42300,
		3080	=>	42303,
		3081	=>	42306,
		3082	=>	42309,
		3083	=>	42312,
		3084	=>	42315,
		3085	=>	42318,
		3086	=>	42321,
		3087	=>	42324,
		3088	=>	42327,
		3089	=>	42330,
		3090	=>	42334,
		3091	=>	42337,
		3092	=>	42340,
		3093	=>	42343,
		3094	=>	42346,
		3095	=>	42349,
		3096	=>	42352,
		3097	=>	42355,
		3098	=>	42358,
		3099	=>	42361,
		3100	=>	42364,
		3101	=>	42367,
		3102	=>	42370,
		3103	=>	42373,
		3104	=>	42376,
		3105	=>	42379,
		3106	=>	42382,
		3107	=>	42385,
		3108	=>	42388,
		3109	=>	42391,
		3110	=>	42394,
		3111	=>	42397,
		3112	=>	42400,
		3113	=>	42403,
		3114	=>	42406,
		3115	=>	42409,
		3116	=>	42412,
		3117	=>	42415,
		3118	=>	42418,
		3119	=>	42421,
		3120	=>	42424,
		3121	=>	42427,
		3122	=>	42430,
		3123	=>	42433,
		3124	=>	42436,
		3125	=>	42439,
		3126	=>	42442,
		3127	=>	42445,
		3128	=>	42448,
		3129	=>	42451,
		3130	=>	42454,
		3131	=>	42457,
		3132	=>	42460,
		3133	=>	42463,
		3134	=>	42466,
		3135	=>	42469,
		3136	=>	42472,
		3137	=>	42475,
		3138	=>	42478,
		3139	=>	42481,
		3140	=>	42484,
		3141	=>	42487,
		3142	=>	42490,
		3143	=>	42493,
		3144	=>	42496,
		3145	=>	42499,
		3146	=>	42502,
		3147	=>	42505,
		3148	=>	42508,
		3149	=>	42511,
		3150	=>	42514,
		3151	=>	42517,
		3152	=>	42520,
		3153	=>	42523,
		3154	=>	42526,
		3155	=>	42529,
		3156	=>	42532,
		3157	=>	42535,
		3158	=>	42538,
		3159	=>	42541,
		3160	=>	42544,
		3161	=>	42547,
		3162	=>	42550,
		3163	=>	42553,
		3164	=>	42556,
		3165	=>	42559,
		3166	=>	42562,
		3167	=>	42565,
		3168	=>	42568,
		3169	=>	42571,
		3170	=>	42574,
		3171	=>	42577,
		3172	=>	42580,
		3173	=>	42583,
		3174	=>	42586,
		3175	=>	42589,
		3176	=>	42592,
		3177	=>	42595,
		3178	=>	42598,
		3179	=>	42601,
		3180	=>	42604,
		3181	=>	42607,
		3182	=>	42610,
		3183	=>	42613,
		3184	=>	42616,
		3185	=>	42619,
		3186	=>	42622,
		3187	=>	42625,
		3188	=>	42628,
		3189	=>	42631,
		3190	=>	42634,
		3191	=>	42637,
		3192	=>	42640,
		3193	=>	42643,
		3194	=>	42646,
		3195	=>	42649,
		3196	=>	42651,
		3197	=>	42654,
		3198	=>	42657,
		3199	=>	42660,
		3200	=>	42663,
		3201	=>	42666,
		3202	=>	42669,
		3203	=>	42672,
		3204	=>	42675,
		3205	=>	42678,
		3206	=>	42681,
		3207	=>	42684,
		3208	=>	42687,
		3209	=>	42690,
		3210	=>	42693,
		3211	=>	42696,
		3212	=>	42699,
		3213	=>	42702,
		3214	=>	42705,
		3215	=>	42708,
		3216	=>	42711,
		3217	=>	42714,
		3218	=>	42717,
		3219	=>	42720,
		3220	=>	42723,
		3221	=>	42726,
		3222	=>	42729,
		3223	=>	42732,
		3224	=>	42735,
		3225	=>	42738,
		3226	=>	42741,
		3227	=>	42744,
		3228	=>	42747,
		3229	=>	42750,
		3230	=>	42753,
		3231	=>	42756,
		3232	=>	42759,
		3233	=>	42762,
		3234	=>	42765,
		3235	=>	42768,
		3236	=>	42771,
		3237	=>	42774,
		3238	=>	42777,
		3239	=>	42780,
		3240	=>	42783,
		3241	=>	42786,
		3242	=>	42789,
		3243	=>	42792,
		3244	=>	42795,
		3245	=>	42798,
		3246	=>	42801,
		3247	=>	42804,
		3248	=>	42807,
		3249	=>	42810,
		3250	=>	42813,
		3251	=>	42816,
		3252	=>	42819,
		3253	=>	42822,
		3254	=>	42825,
		3255	=>	42828,
		3256	=>	42831,
		3257	=>	42834,
		3258	=>	42837,
		3259	=>	42840,
		3260	=>	42843,
		3261	=>	42846,
		3262	=>	42849,
		3263	=>	42852,
		3264	=>	42855,
		3265	=>	42858,
		3266	=>	42861,
		3267	=>	42864,
		3268	=>	42867,
		3269	=>	42870,
		3270	=>	42873,
		3271	=>	42876,
		3272	=>	42879,
		3273	=>	42882,
		3274	=>	42885,
		3275	=>	42888,
		3276	=>	42891,
		3277	=>	42894,
		3278	=>	42897,
		3279	=>	42900,
		3280	=>	42903,
		3281	=>	42906,
		3282	=>	42909,
		3283	=>	42912,
		3284	=>	42915,
		3285	=>	42918,
		3286	=>	42921,
		3287	=>	42924,
		3288	=>	42927,
		3289	=>	42930,
		3290	=>	42933,
		3291	=>	42936,
		3292	=>	42939,
		3293	=>	42942,
		3294	=>	42945,
		3295	=>	42948,
		3296	=>	42951,
		3297	=>	42954,
		3298	=>	42957,
		3299	=>	42960,
		3300	=>	42963,
		3301	=>	42965,
		3302	=>	42968,
		3303	=>	42971,
		3304	=>	42974,
		3305	=>	42977,
		3306	=>	42980,
		3307	=>	42983,
		3308	=>	42986,
		3309	=>	42989,
		3310	=>	42992,
		3311	=>	42995,
		3312	=>	42998,
		3313	=>	43001,
		3314	=>	43004,
		3315	=>	43007,
		3316	=>	43010,
		3317	=>	43013,
		3318	=>	43016,
		3319	=>	43019,
		3320	=>	43022,
		3321	=>	43025,
		3322	=>	43028,
		3323	=>	43031,
		3324	=>	43034,
		3325	=>	43037,
		3326	=>	43040,
		3327	=>	43043,
		3328	=>	43046,
		3329	=>	43049,
		3330	=>	43052,
		3331	=>	43055,
		3332	=>	43058,
		3333	=>	43061,
		3334	=>	43064,
		3335	=>	43067,
		3336	=>	43070,
		3337	=>	43073,
		3338	=>	43076,
		3339	=>	43079,
		3340	=>	43082,
		3341	=>	43085,
		3342	=>	43088,
		3343	=>	43091,
		3344	=>	43094,
		3345	=>	43097,
		3346	=>	43100,
		3347	=>	43103,
		3348	=>	43106,
		3349	=>	43109,
		3350	=>	43112,
		3351	=>	43115,
		3352	=>	43118,
		3353	=>	43121,
		3354	=>	43124,
		3355	=>	43127,
		3356	=>	43130,
		3357	=>	43133,
		3358	=>	43136,
		3359	=>	43138,
		3360	=>	43141,
		3361	=>	43144,
		3362	=>	43147,
		3363	=>	43150,
		3364	=>	43153,
		3365	=>	43156,
		3366	=>	43159,
		3367	=>	43162,
		3368	=>	43165,
		3369	=>	43168,
		3370	=>	43171,
		3371	=>	43174,
		3372	=>	43177,
		3373	=>	43180,
		3374	=>	43183,
		3375	=>	43186,
		3376	=>	43189,
		3377	=>	43192,
		3378	=>	43195,
		3379	=>	43198,
		3380	=>	43201,
		3381	=>	43204,
		3382	=>	43207,
		3383	=>	43210,
		3384	=>	43213,
		3385	=>	43216,
		3386	=>	43219,
		3387	=>	43222,
		3388	=>	43225,
		3389	=>	43228,
		3390	=>	43231,
		3391	=>	43234,
		3392	=>	43237,
		3393	=>	43240,
		3394	=>	43243,
		3395	=>	43246,
		3396	=>	43249,
		3397	=>	43252,
		3398	=>	43255,
		3399	=>	43258,
		3400	=>	43261,
		3401	=>	43264,
		3402	=>	43267,
		3403	=>	43270,
		3404	=>	43272,
		3405	=>	43275,
		3406	=>	43278,
		3407	=>	43281,
		3408	=>	43284,
		3409	=>	43287,
		3410	=>	43290,
		3411	=>	43293,
		3412	=>	43296,
		3413	=>	43299,
		3414	=>	43302,
		3415	=>	43305,
		3416	=>	43308,
		3417	=>	43311,
		3418	=>	43314,
		3419	=>	43317,
		3420	=>	43320,
		3421	=>	43323,
		3422	=>	43326,
		3423	=>	43329,
		3424	=>	43332,
		3425	=>	43335,
		3426	=>	43338,
		3427	=>	43341,
		3428	=>	43344,
		3429	=>	43347,
		3430	=>	43350,
		3431	=>	43353,
		3432	=>	43356,
		3433	=>	43359,
		3434	=>	43362,
		3435	=>	43365,
		3436	=>	43368,
		3437	=>	43371,
		3438	=>	43374,
		3439	=>	43377,
		3440	=>	43380,
		3441	=>	43383,
		3442	=>	43386,
		3443	=>	43388,
		3444	=>	43391,
		3445	=>	43394,
		3446	=>	43397,
		3447	=>	43400,
		3448	=>	43403,
		3449	=>	43406,
		3450	=>	43409,
		3451	=>	43412,
		3452	=>	43415,
		3453	=>	43418,
		3454	=>	43421,
		3455	=>	43424,
		3456	=>	43427,
		3457	=>	43430,
		3458	=>	43433,
		3459	=>	43436,
		3460	=>	43439,
		3461	=>	43442,
		3462	=>	43445,
		3463	=>	43448,
		3464	=>	43451,
		3465	=>	43454,
		3466	=>	43457,
		3467	=>	43460,
		3468	=>	43463,
		3469	=>	43466,
		3470	=>	43469,
		3471	=>	43472,
		3472	=>	43475,
		3473	=>	43478,
		3474	=>	43481,
		3475	=>	43484,
		3476	=>	43486,
		3477	=>	43489,
		3478	=>	43492,
		3479	=>	43495,
		3480	=>	43498,
		3481	=>	43501,
		3482	=>	43504,
		3483	=>	43507,
		3484	=>	43510,
		3485	=>	43513,
		3486	=>	43516,
		3487	=>	43519,
		3488	=>	43522,
		3489	=>	43525,
		3490	=>	43528,
		3491	=>	43531,
		3492	=>	43534,
		3493	=>	43537,
		3494	=>	43540,
		3495	=>	43543,
		3496	=>	43546,
		3497	=>	43549,
		3498	=>	43552,
		3499	=>	43555,
		3500	=>	43558,
		3501	=>	43561,
		3502	=>	43564,
		3503	=>	43567,
		3504	=>	43570,
		3505	=>	43573,
		3506	=>	43576,
		3507	=>	43578,
		3508	=>	43581,
		3509	=>	43584,
		3510	=>	43587,
		3511	=>	43590,
		3512	=>	43593,
		3513	=>	43596,
		3514	=>	43599,
		3515	=>	43602,
		3516	=>	43605,
		3517	=>	43608,
		3518	=>	43611,
		3519	=>	43614,
		3520	=>	43617,
		3521	=>	43620,
		3522	=>	43623,
		3523	=>	43626,
		3524	=>	43629,
		3525	=>	43632,
		3526	=>	43635,
		3527	=>	43638,
		3528	=>	43641,
		3529	=>	43644,
		3530	=>	43647,
		3531	=>	43650,
		3532	=>	43653,
		3533	=>	43656,
		3534	=>	43659,
		3535	=>	43661,
		3536	=>	43664,
		3537	=>	43667,
		3538	=>	43670,
		3539	=>	43673,
		3540	=>	43676,
		3541	=>	43679,
		3542	=>	43682,
		3543	=>	43685,
		3544	=>	43688,
		3545	=>	43691,
		3546	=>	43694,
		3547	=>	43697,
		3548	=>	43700,
		3549	=>	43703,
		3550	=>	43706,
		3551	=>	43709,
		3552	=>	43712,
		3553	=>	43715,
		3554	=>	43718,
		3555	=>	43721,
		3556	=>	43724,
		3557	=>	43727,
		3558	=>	43730,
		3559	=>	43733,
		3560	=>	43736,
		3561	=>	43738,
		3562	=>	43741,
		3563	=>	43744,
		3564	=>	43747,
		3565	=>	43750,
		3566	=>	43753,
		3567	=>	43756,
		3568	=>	43759,
		3569	=>	43762,
		3570	=>	43765,
		3571	=>	43768,
		3572	=>	43771,
		3573	=>	43774,
		3574	=>	43777,
		3575	=>	43780,
		3576	=>	43783,
		3577	=>	43786,
		3578	=>	43789,
		3579	=>	43792,
		3580	=>	43795,
		3581	=>	43798,
		3582	=>	43801,
		3583	=>	43804,
		3584	=>	43807,
		3585	=>	43809,
		3586	=>	43812,
		3587	=>	43815,
		3588	=>	43818,
		3589	=>	43821,
		3590	=>	43824,
		3591	=>	43827,
		3592	=>	43830,
		3593	=>	43833,
		3594	=>	43836,
		3595	=>	43839,
		3596	=>	43842,
		3597	=>	43845,
		3598	=>	43848,
		3599	=>	43851,
		3600	=>	43854,
		3601	=>	43857,
		3602	=>	43860,
		3603	=>	43863,
		3604	=>	43866,
		3605	=>	43869,
		3606	=>	43872,
		3607	=>	43875,
		3608	=>	43877,
		3609	=>	43880,
		3610	=>	43883,
		3611	=>	43886,
		3612	=>	43889,
		3613	=>	43892,
		3614	=>	43895,
		3615	=>	43898,
		3616	=>	43901,
		3617	=>	43904,
		3618	=>	43907,
		3619	=>	43910,
		3620	=>	43913,
		3621	=>	43916,
		3622	=>	43919,
		3623	=>	43922,
		3624	=>	43925,
		3625	=>	43928,
		3626	=>	43931,
		3627	=>	43934,
		3628	=>	43937,
		3629	=>	43940,
		3630	=>	43942,
		3631	=>	43945,
		3632	=>	43948,
		3633	=>	43951,
		3634	=>	43954,
		3635	=>	43957,
		3636	=>	43960,
		3637	=>	43963,
		3638	=>	43966,
		3639	=>	43969,
		3640	=>	43972,
		3641	=>	43975,
		3642	=>	43978,
		3643	=>	43981,
		3644	=>	43984,
		3645	=>	43987,
		3646	=>	43990,
		3647	=>	43993,
		3648	=>	43996,
		3649	=>	43999,
		3650	=>	44002,
		3651	=>	44004,
		3652	=>	44007,
		3653	=>	44010,
		3654	=>	44013,
		3655	=>	44016,
		3656	=>	44019,
		3657	=>	44022,
		3658	=>	44025,
		3659	=>	44028,
		3660	=>	44031,
		3661	=>	44034,
		3662	=>	44037,
		3663	=>	44040,
		3664	=>	44043,
		3665	=>	44046,
		3666	=>	44049,
		3667	=>	44052,
		3668	=>	44055,
		3669	=>	44058,
		3670	=>	44061,
		3671	=>	44063,
		3672	=>	44066,
		3673	=>	44069,
		3674	=>	44072,
		3675	=>	44075,
		3676	=>	44078,
		3677	=>	44081,
		3678	=>	44084,
		3679	=>	44087,
		3680	=>	44090,
		3681	=>	44093,
		3682	=>	44096,
		3683	=>	44099,
		3684	=>	44102,
		3685	=>	44105,
		3686	=>	44108,
		3687	=>	44111,
		3688	=>	44114,
		3689	=>	44117,
		3690	=>	44120,
		3691	=>	44122,
		3692	=>	44125,
		3693	=>	44128,
		3694	=>	44131,
		3695	=>	44134,
		3696	=>	44137,
		3697	=>	44140,
		3698	=>	44143,
		3699	=>	44146,
		3700	=>	44149,
		3701	=>	44152,
		3702	=>	44155,
		3703	=>	44158,
		3704	=>	44161,
		3705	=>	44164,
		3706	=>	44167,
		3707	=>	44170,
		3708	=>	44173,
		3709	=>	44175,
		3710	=>	44178,
		3711	=>	44181,
		3712	=>	44184,
		3713	=>	44187,
		3714	=>	44190,
		3715	=>	44193,
		3716	=>	44196,
		3717	=>	44199,
		3718	=>	44202,
		3719	=>	44205,
		3720	=>	44208,
		3721	=>	44211,
		3722	=>	44214,
		3723	=>	44217,
		3724	=>	44220,
		3725	=>	44223,
		3726	=>	44226,
		3727	=>	44228,
		3728	=>	44231,
		3729	=>	44234,
		3730	=>	44237,
		3731	=>	44240,
		3732	=>	44243,
		3733	=>	44246,
		3734	=>	44249,
		3735	=>	44252,
		3736	=>	44255,
		3737	=>	44258,
		3738	=>	44261,
		3739	=>	44264,
		3740	=>	44267,
		3741	=>	44270,
		3742	=>	44273,
		3743	=>	44276,
		3744	=>	44278,
		3745	=>	44281,
		3746	=>	44284,
		3747	=>	44287,
		3748	=>	44290,
		3749	=>	44293,
		3750	=>	44296,
		3751	=>	44299,
		3752	=>	44302,
		3753	=>	44305,
		3754	=>	44308,
		3755	=>	44311,
		3756	=>	44314,
		3757	=>	44317,
		3758	=>	44320,
		3759	=>	44323,
		3760	=>	44326,
		3761	=>	44328,
		3762	=>	44331,
		3763	=>	44334,
		3764	=>	44337,
		3765	=>	44340,
		3766	=>	44343,
		3767	=>	44346,
		3768	=>	44349,
		3769	=>	44352,
		3770	=>	44355,
		3771	=>	44358,
		3772	=>	44361,
		3773	=>	44364,
		3774	=>	44367,
		3775	=>	44370,
		3776	=>	44373,
		3777	=>	44375,
		3778	=>	44378,
		3779	=>	44381,
		3780	=>	44384,
		3781	=>	44387,
		3782	=>	44390,
		3783	=>	44393,
		3784	=>	44396,
		3785	=>	44399,
		3786	=>	44402,
		3787	=>	44405,
		3788	=>	44408,
		3789	=>	44411,
		3790	=>	44414,
		3791	=>	44417,
		3792	=>	44420,
		3793	=>	44422,
		3794	=>	44425,
		3795	=>	44428,
		3796	=>	44431,
		3797	=>	44434,
		3798	=>	44437,
		3799	=>	44440,
		3800	=>	44443,
		3801	=>	44446,
		3802	=>	44449,
		3803	=>	44452,
		3804	=>	44455,
		3805	=>	44458,
		3806	=>	44461,
		3807	=>	44464,
		3808	=>	44467,
		3809	=>	44469,
		3810	=>	44472,
		3811	=>	44475,
		3812	=>	44478,
		3813	=>	44481,
		3814	=>	44484,
		3815	=>	44487,
		3816	=>	44490,
		3817	=>	44493,
		3818	=>	44496,
		3819	=>	44499,
		3820	=>	44502,
		3821	=>	44505,
		3822	=>	44508,
		3823	=>	44511,
		3824	=>	44513,
		3825	=>	44516,
		3826	=>	44519,
		3827	=>	44522,
		3828	=>	44525,
		3829	=>	44528,
		3830	=>	44531,
		3831	=>	44534,
		3832	=>	44537,
		3833	=>	44540,
		3834	=>	44543,
		3835	=>	44546,
		3836	=>	44549,
		3837	=>	44552,
		3838	=>	44554,
		3839	=>	44557,
		3840	=>	44560,
		3841	=>	44563,
		3842	=>	44566,
		3843	=>	44569,
		3844	=>	44572,
		3845	=>	44575,
		3846	=>	44578,
		3847	=>	44581,
		3848	=>	44584,
		3849	=>	44587,
		3850	=>	44590,
		3851	=>	44593,
		3852	=>	44596,
		3853	=>	44598,
		3854	=>	44601,
		3855	=>	44604,
		3856	=>	44607,
		3857	=>	44610,
		3858	=>	44613,
		3859	=>	44616,
		3860	=>	44619,
		3861	=>	44622,
		3862	=>	44625,
		3863	=>	44628,
		3864	=>	44631,
		3865	=>	44634,
		3866	=>	44637,
		3867	=>	44639,
		3868	=>	44642,
		3869	=>	44645,
		3870	=>	44648,
		3871	=>	44651,
		3872	=>	44654,
		3873	=>	44657,
		3874	=>	44660,
		3875	=>	44663,
		3876	=>	44666,
		3877	=>	44669,
		3878	=>	44672,
		3879	=>	44675,
		3880	=>	44678,
		3881	=>	44680,
		3882	=>	44683,
		3883	=>	44686,
		3884	=>	44689,
		3885	=>	44692,
		3886	=>	44695,
		3887	=>	44698,
		3888	=>	44701,
		3889	=>	44704,
		3890	=>	44707,
		3891	=>	44710,
		3892	=>	44713,
		3893	=>	44716,
		3894	=>	44718,
		3895	=>	44721,
		3896	=>	44724,
		3897	=>	44727,
		3898	=>	44730,
		3899	=>	44733,
		3900	=>	44736,
		3901	=>	44739,
		3902	=>	44742,
		3903	=>	44745,
		3904	=>	44748,
		3905	=>	44751,
		3906	=>	44754,
		3907	=>	44756,
		3908	=>	44759,
		3909	=>	44762,
		3910	=>	44765,
		3911	=>	44768,
		3912	=>	44771,
		3913	=>	44774,
		3914	=>	44777,
		3915	=>	44780,
		3916	=>	44783,
		3917	=>	44786,
		3918	=>	44789,
		3919	=>	44792,
		3920	=>	44794,
		3921	=>	44797,
		3922	=>	44800,
		3923	=>	44803,
		3924	=>	44806,
		3925	=>	44809,
		3926	=>	44812,
		3927	=>	44815,
		3928	=>	44818,
		3929	=>	44821,
		3930	=>	44824,
		3931	=>	44827,
		3932	=>	44830,
		3933	=>	44832,
		3934	=>	44835,
		3935	=>	44838,
		3936	=>	44841,
		3937	=>	44844,
		3938	=>	44847,
		3939	=>	44850,
		3940	=>	44853,
		3941	=>	44856,
		3942	=>	44859,
		3943	=>	44862,
		3944	=>	44865,
		3945	=>	44868,
		3946	=>	44870,
		3947	=>	44873,
		3948	=>	44876,
		3949	=>	44879,
		3950	=>	44882,
		3951	=>	44885,
		3952	=>	44888,
		3953	=>	44891,
		3954	=>	44894,
		3955	=>	44897,
		3956	=>	44900,
		3957	=>	44903,
		3958	=>	44905,
		3959	=>	44908,
		3960	=>	44911,
		3961	=>	44914,
		3962	=>	44917,
		3963	=>	44920,
		3964	=>	44923,
		3965	=>	44926,
		3966	=>	44929,
		3967	=>	44932,
		3968	=>	44935,
		3969	=>	44938,
		3970	=>	44940,
		3971	=>	44943,
		3972	=>	44946,
		3973	=>	44949,
		3974	=>	44952,
		3975	=>	44955,
		3976	=>	44958,
		3977	=>	44961,
		3978	=>	44964,
		3979	=>	44967,
		3980	=>	44970,
		3981	=>	44973,
		3982	=>	44975,
		3983	=>	44978,
		3984	=>	44981,
		3985	=>	44984,
		3986	=>	44987,
		3987	=>	44990,
		3988	=>	44993,
		3989	=>	44996,
		3990	=>	44999,
		3991	=>	45002,
		3992	=>	45005,
		3993	=>	45008,
		3994	=>	45010,
		3995	=>	45013,
		3996	=>	45016,
		3997	=>	45019,
		3998	=>	45022,
		3999	=>	45025,
		4000	=>	45028,
		4001	=>	45031,
		4002	=>	45034,
		4003	=>	45037,
		4004	=>	45040,
		4005	=>	45042,
		4006	=>	45045,
		4007	=>	45048,
		4008	=>	45051,
		4009	=>	45054,
		4010	=>	45057,
		4011	=>	45060,
		4012	=>	45063,
		4013	=>	45066,
		4014	=>	45069,
		4015	=>	45072,
		4016	=>	45075,
		4017	=>	45077,
		4018	=>	45080,
		4019	=>	45083,
		4020	=>	45086,
		4021	=>	45089,
		4022	=>	45092,
		4023	=>	45095,
		4024	=>	45098,
		4025	=>	45101,
		4026	=>	45104,
		4027	=>	45107,
		4028	=>	45109,
		4029	=>	45112,
		4030	=>	45115,
		4031	=>	45118,
		4032	=>	45121,
		4033	=>	45124,
		4034	=>	45127,
		4035	=>	45130,
		4036	=>	45133,
		4037	=>	45136,
		4038	=>	45139,
		4039	=>	45141,
		4040	=>	45144,
		4041	=>	45147,
		4042	=>	45150,
		4043	=>	45153,
		4044	=>	45156,
		4045	=>	45159,
		4046	=>	45162,
		4047	=>	45165,
		4048	=>	45168,
		4049	=>	45171,
		4050	=>	45173,
		4051	=>	45176,
		4052	=>	45179,
		4053	=>	45182,
		4054	=>	45185,
		4055	=>	45188,
		4056	=>	45191,
		4057	=>	45194,
		4058	=>	45197,
		4059	=>	45200,
		4060	=>	45203,
		4061	=>	45205,
		4062	=>	45208,
		4063	=>	45211,
		4064	=>	45214,
		4065	=>	45217,
		4066	=>	45220,
		4067	=>	45223,
		4068	=>	45226,
		4069	=>	45229,
		4070	=>	45232,
		4071	=>	45234,
		4072	=>	45237,
		4073	=>	45240,
		4074	=>	45243,
		4075	=>	45246,
		4076	=>	45249,
		4077	=>	45252,
		4078	=>	45255,
		4079	=>	45258,
		4080	=>	45261,
		4081	=>	45264,
		4082	=>	45266,
		4083	=>	45269,
		4084	=>	45272,
		4085	=>	45275,
		4086	=>	45278,
		4087	=>	45281,
		4088	=>	45284,
		4089	=>	45287,
		4090	=>	45290,
		4091	=>	45293,
		4092	=>	45295,
		4093	=>	45298,
		4094	=>	45301,
		4095	=>	45304,
		4096	=>	45307,
		4097	=>	45310,
		4098	=>	45313,
		4099	=>	45316,
		4100	=>	45319,
		4101	=>	45322,
		4102	=>	45324,
		4103	=>	45327,
		4104	=>	45330,
		4105	=>	45333,
		4106	=>	45336,
		4107	=>	45339,
		4108	=>	45342,
		4109	=>	45345,
		4110	=>	45348,
		4111	=>	45351,
		4112	=>	45354,
		4113	=>	45356,
		4114	=>	45359,
		4115	=>	45362,
		4116	=>	45365,
		4117	=>	45368,
		4118	=>	45371,
		4119	=>	45374,
		4120	=>	45377,
		4121	=>	45380,
		4122	=>	45383,
		4123	=>	45385,
		4124	=>	45388,
		4125	=>	45391,
		4126	=>	45394,
		4127	=>	45397,
		4128	=>	45400,
		4129	=>	45403,
		4130	=>	45406,
		4131	=>	45409,
		4132	=>	45411,
		4133	=>	45414,
		4134	=>	45417,
		4135	=>	45420,
		4136	=>	45423,
		4137	=>	45426,
		4138	=>	45429,
		4139	=>	45432,
		4140	=>	45435,
		4141	=>	45438,
		4142	=>	45440,
		4143	=>	45443,
		4144	=>	45446,
		4145	=>	45449,
		4146	=>	45452,
		4147	=>	45455,
		4148	=>	45458,
		4149	=>	45461,
		4150	=>	45464,
		4151	=>	45467,
		4152	=>	45469,
		4153	=>	45472,
		4154	=>	45475,
		4155	=>	45478,
		4156	=>	45481,
		4157	=>	45484,
		4158	=>	45487,
		4159	=>	45490,
		4160	=>	45493,
		4161	=>	45495,
		4162	=>	45498,
		4163	=>	45501,
		4164	=>	45504,
		4165	=>	45507,
		4166	=>	45510,
		4167	=>	45513,
		4168	=>	45516,
		4169	=>	45519,
		4170	=>	45522,
		4171	=>	45524,
		4172	=>	45527,
		4173	=>	45530,
		4174	=>	45533,
		4175	=>	45536,
		4176	=>	45539,
		4177	=>	45542,
		4178	=>	45545,
		4179	=>	45548,
		4180	=>	45550,
		4181	=>	45553,
		4182	=>	45556,
		4183	=>	45559,
		4184	=>	45562,
		4185	=>	45565,
		4186	=>	45568,
		4187	=>	45571,
		4188	=>	45574,
		4189	=>	45577,
		4190	=>	45579,
		4191	=>	45582,
		4192	=>	45585,
		4193	=>	45588,
		4194	=>	45591,
		4195	=>	45594,
		4196	=>	45597,
		4197	=>	45600,
		4198	=>	45603,
		4199	=>	45605,
		4200	=>	45608,
		4201	=>	45611,
		4202	=>	45614,
		4203	=>	45617,
		4204	=>	45620,
		4205	=>	45623,
		4206	=>	45626,
		4207	=>	45629,
		4208	=>	45631,
		4209	=>	45634,
		4210	=>	45637,
		4211	=>	45640,
		4212	=>	45643,
		4213	=>	45646,
		4214	=>	45649,
		4215	=>	45652,
		4216	=>	45655,
		4217	=>	45657,
		4218	=>	45660,
		4219	=>	45663,
		4220	=>	45666,
		4221	=>	45669,
		4222	=>	45672,
		4223	=>	45675,
		4224	=>	45678,
		4225	=>	45681,
		4226	=>	45683,
		4227	=>	45686,
		4228	=>	45689,
		4229	=>	45692,
		4230	=>	45695,
		4231	=>	45698,
		4232	=>	45701,
		4233	=>	45704,
		4234	=>	45707,
		4235	=>	45709,
		4236	=>	45712,
		4237	=>	45715,
		4238	=>	45718,
		4239	=>	45721,
		4240	=>	45724,
		4241	=>	45727,
		4242	=>	45730,
		4243	=>	45732,
		4244	=>	45735,
		4245	=>	45738,
		4246	=>	45741,
		4247	=>	45744,
		4248	=>	45747,
		4249	=>	45750,
		4250	=>	45753,
		4251	=>	45756,
		4252	=>	45758,
		4253	=>	45761,
		4254	=>	45764,
		4255	=>	45767,
		4256	=>	45770,
		4257	=>	45773,
		4258	=>	45776,
		4259	=>	45779,
		4260	=>	45782,
		4261	=>	45784,
		4262	=>	45787,
		4263	=>	45790,
		4264	=>	45793,
		4265	=>	45796,
		4266	=>	45799,
		4267	=>	45802,
		4268	=>	45805,
		4269	=>	45807,
		4270	=>	45810,
		4271	=>	45813,
		4272	=>	45816,
		4273	=>	45819,
		4274	=>	45822,
		4275	=>	45825,
		4276	=>	45828,
		4277	=>	45831,
		4278	=>	45833,
		4279	=>	45836,
		4280	=>	45839,
		4281	=>	45842,
		4282	=>	45845,
		4283	=>	45848,
		4284	=>	45851,
		4285	=>	45854,
		4286	=>	45856,
		4287	=>	45859,
		4288	=>	45862,
		4289	=>	45865,
		4290	=>	45868,
		4291	=>	45871,
		4292	=>	45874,
		4293	=>	45877,
		4294	=>	45879,
		4295	=>	45882,
		4296	=>	45885,
		4297	=>	45888,
		4298	=>	45891,
		4299	=>	45894,
		4300	=>	45897,
		4301	=>	45900,
		4302	=>	45902,
		4303	=>	45905,
		4304	=>	45908,
		4305	=>	45911,
		4306	=>	45914,
		4307	=>	45917,
		4308	=>	45920,
		4309	=>	45923,
		4310	=>	45926,
		4311	=>	45928,
		4312	=>	45931,
		4313	=>	45934,
		4314	=>	45937,
		4315	=>	45940,
		4316	=>	45943,
		4317	=>	45946,
		4318	=>	45949,
		4319	=>	45951,
		4320	=>	45954,
		4321	=>	45957,
		4322	=>	45960,
		4323	=>	45963,
		4324	=>	45966,
		4325	=>	45969,
		4326	=>	45972,
		4327	=>	45974,
		4328	=>	45977,
		4329	=>	45980,
		4330	=>	45983,
		4331	=>	45986,
		4332	=>	45989,
		4333	=>	45992,
		4334	=>	45995,
		4335	=>	45997,
		4336	=>	46000,
		4337	=>	46003,
		4338	=>	46006,
		4339	=>	46009,
		4340	=>	46012,
		4341	=>	46015,
		4342	=>	46018,
		4343	=>	46020,
		4344	=>	46023,
		4345	=>	46026,
		4346	=>	46029,
		4347	=>	46032,
		4348	=>	46035,
		4349	=>	46038,
		4350	=>	46041,
		4351	=>	46043,
		4352	=>	46046,
		4353	=>	46049,
		4354	=>	46052,
		4355	=>	46055,
		4356	=>	46058,
		4357	=>	46061,
		4358	=>	46063,
		4359	=>	46066,
		4360	=>	46069,
		4361	=>	46072,
		4362	=>	46075,
		4363	=>	46078,
		4364	=>	46081,
		4365	=>	46084,
		4366	=>	46086,
		4367	=>	46089,
		4368	=>	46092,
		4369	=>	46095,
		4370	=>	46098,
		4371	=>	46101,
		4372	=>	46104,
		4373	=>	46107,
		4374	=>	46109,
		4375	=>	46112,
		4376	=>	46115,
		4377	=>	46118,
		4378	=>	46121,
		4379	=>	46124,
		4380	=>	46127,
		4381	=>	46129,
		4382	=>	46132,
		4383	=>	46135,
		4384	=>	46138,
		4385	=>	46141,
		4386	=>	46144,
		4387	=>	46147,
		4388	=>	46150,
		4389	=>	46152,
		4390	=>	46155,
		4391	=>	46158,
		4392	=>	46161,
		4393	=>	46164,
		4394	=>	46167,
		4395	=>	46170,
		4396	=>	46172,
		4397	=>	46175,
		4398	=>	46178,
		4399	=>	46181,
		4400	=>	46184,
		4401	=>	46187,
		4402	=>	46190,
		4403	=>	46193,
		4404	=>	46195,
		4405	=>	46198,
		4406	=>	46201,
		4407	=>	46204,
		4408	=>	46207,
		4409	=>	46210,
		4410	=>	46213,
		4411	=>	46215,
		4412	=>	46218,
		4413	=>	46221,
		4414	=>	46224,
		4415	=>	46227,
		4416	=>	46230,
		4417	=>	46233,
		4418	=>	46236,
		4419	=>	46238,
		4420	=>	46241,
		4421	=>	46244,
		4422	=>	46247,
		4423	=>	46250,
		4424	=>	46253,
		4425	=>	46256,
		4426	=>	46258,
		4427	=>	46261,
		4428	=>	46264,
		4429	=>	46267,
		4430	=>	46270,
		4431	=>	46273,
		4432	=>	46276,
		4433	=>	46278,
		4434	=>	46281,
		4435	=>	46284,
		4436	=>	46287,
		4437	=>	46290,
		4438	=>	46293,
		4439	=>	46296,
		4440	=>	46299,
		4441	=>	46301,
		4442	=>	46304,
		4443	=>	46307,
		4444	=>	46310,
		4445	=>	46313,
		4446	=>	46316,
		4447	=>	46319,
		4448	=>	46321,
		4449	=>	46324,
		4450	=>	46327,
		4451	=>	46330,
		4452	=>	46333,
		4453	=>	46336,
		4454	=>	46339,
		4455	=>	46341,
		4456	=>	46344,
		4457	=>	46347,
		4458	=>	46350,
		4459	=>	46353,
		4460	=>	46356,
		4461	=>	46359,
		4462	=>	46361,
		4463	=>	46364,
		4464	=>	46367,
		4465	=>	46370,
		4466	=>	46373,
		4467	=>	46376,
		4468	=>	46379,
		4469	=>	46381,
		4470	=>	46384,
		4471	=>	46387,
		4472	=>	46390,
		4473	=>	46393,
		4474	=>	46396,
		4475	=>	46399,
		4476	=>	46401,
		4477	=>	46404,
		4478	=>	46407,
		4479	=>	46410,
		4480	=>	46413,
		4481	=>	46416,
		4482	=>	46419,
		4483	=>	46421,
		4484	=>	46424,
		4485	=>	46427,
		4486	=>	46430,
		4487	=>	46433,
		4488	=>	46436,
		4489	=>	46439,
		4490	=>	46441,
		4491	=>	46444,
		4492	=>	46447,
		4493	=>	46450,
		4494	=>	46453,
		4495	=>	46456,
		4496	=>	46459,
		4497	=>	46461,
		4498	=>	46464,
		4499	=>	46467,
		4500	=>	46470,
		4501	=>	46473,
		4502	=>	46476,
		4503	=>	46479,
		4504	=>	46481,
		4505	=>	46484,
		4506	=>	46487,
		4507	=>	46490,
		4508	=>	46493,
		4509	=>	46496,
		4510	=>	46498,
		4511	=>	46501,
		4512	=>	46504,
		4513	=>	46507,
		4514	=>	46510,
		4515	=>	46513,
		4516	=>	46516,
		4517	=>	46518,
		4518	=>	46521,
		4519	=>	46524,
		4520	=>	46527,
		4521	=>	46530,
		4522	=>	46533,
		4523	=>	46536,
		4524	=>	46538,
		4525	=>	46541,
		4526	=>	46544,
		4527	=>	46547,
		4528	=>	46550,
		4529	=>	46553,
		4530	=>	46556,
		4531	=>	46558,
		4532	=>	46561,
		4533	=>	46564,
		4534	=>	46567,
		4535	=>	46570,
		4536	=>	46573,
		4537	=>	46575,
		4538	=>	46578,
		4539	=>	46581,
		4540	=>	46584,
		4541	=>	46587,
		4542	=>	46590,
		4543	=>	46593,
		4544	=>	46595,
		4545	=>	46598,
		4546	=>	46601,
		4547	=>	46604,
		4548	=>	46607,
		4549	=>	46610,
		4550	=>	46612,
		4551	=>	46615,
		4552	=>	46618,
		4553	=>	46621,
		4554	=>	46624,
		4555	=>	46627,
		4556	=>	46630,
		4557	=>	46632,
		4558	=>	46635,
		4559	=>	46638,
		4560	=>	46641,
		4561	=>	46644,
		4562	=>	46647,
		4563	=>	46649,
		4564	=>	46652,
		4565	=>	46655,
		4566	=>	46658,
		4567	=>	46661,
		4568	=>	46664,
		4569	=>	46667,
		4570	=>	46669,
		4571	=>	46672,
		4572	=>	46675,
		4573	=>	46678,
		4574	=>	46681,
		4575	=>	46684,
		4576	=>	46686,
		4577	=>	46689,
		4578	=>	46692,
		4579	=>	46695,
		4580	=>	46698,
		4581	=>	46701,
		4582	=>	46704,
		4583	=>	46706,
		4584	=>	46709,
		4585	=>	46712,
		4586	=>	46715,
		4587	=>	46718,
		4588	=>	46721,
		4589	=>	46723,
		4590	=>	46726,
		4591	=>	46729,
		4592	=>	46732,
		4593	=>	46735,
		4594	=>	46738,
		4595	=>	46740,
		4596	=>	46743,
		4597	=>	46746,
		4598	=>	46749,
		4599	=>	46752,
		4600	=>	46755,
		4601	=>	46758,
		4602	=>	46760,
		4603	=>	46763,
		4604	=>	46766,
		4605	=>	46769,
		4606	=>	46772,
		4607	=>	46775,
		4608	=>	46777,
		4609	=>	46780,
		4610	=>	46783,
		4611	=>	46786,
		4612	=>	46789,
		4613	=>	46792,
		4614	=>	46794,
		4615	=>	46797,
		4616	=>	46800,
		4617	=>	46803,
		4618	=>	46806,
		4619	=>	46809,
		4620	=>	46811,
		4621	=>	46814,
		4622	=>	46817,
		4623	=>	46820,
		4624	=>	46823,
		4625	=>	46826,
		4626	=>	46829,
		4627	=>	46831,
		4628	=>	46834,
		4629	=>	46837,
		4630	=>	46840,
		4631	=>	46843,
		4632	=>	46846,
		4633	=>	46848,
		4634	=>	46851,
		4635	=>	46854,
		4636	=>	46857,
		4637	=>	46860,
		4638	=>	46863,
		4639	=>	46865,
		4640	=>	46868,
		4641	=>	46871,
		4642	=>	46874,
		4643	=>	46877,
		4644	=>	46880,
		4645	=>	46882,
		4646	=>	46885,
		4647	=>	46888,
		4648	=>	46891,
		4649	=>	46894,
		4650	=>	46897,
		4651	=>	46899,
		4652	=>	46902,
		4653	=>	46905,
		4654	=>	46908,
		4655	=>	46911,
		4656	=>	46914,
		4657	=>	46916,
		4658	=>	46919,
		4659	=>	46922,
		4660	=>	46925,
		4661	=>	46928,
		4662	=>	46931,
		4663	=>	46933,
		4664	=>	46936,
		4665	=>	46939,
		4666	=>	46942,
		4667	=>	46945,
		4668	=>	46948,
		4669	=>	46950,
		4670	=>	46953,
		4671	=>	46956,
		4672	=>	46959,
		4673	=>	46962,
		4674	=>	46965,
		4675	=>	46967,
		4676	=>	46970,
		4677	=>	46973,
		4678	=>	46976,
		4679	=>	46979,
		4680	=>	46982,
		4681	=>	46984,
		4682	=>	46987,
		4683	=>	46990,
		4684	=>	46993,
		4685	=>	46996,
		4686	=>	46999,
		4687	=>	47001,
		4688	=>	47004,
		4689	=>	47007,
		4690	=>	47010,
		4691	=>	47013,
		4692	=>	47016,
		4693	=>	47018,
		4694	=>	47021,
		4695	=>	47024,
		4696	=>	47027,
		4697	=>	47030,
		4698	=>	47032,
		4699	=>	47035,
		4700	=>	47038,
		4701	=>	47041,
		4702	=>	47044,
		4703	=>	47047,
		4704	=>	47049,
		4705	=>	47052,
		4706	=>	47055,
		4707	=>	47058,
		4708	=>	47061,
		4709	=>	47064,
		4710	=>	47066,
		4711	=>	47069,
		4712	=>	47072,
		4713	=>	47075,
		4714	=>	47078,
		4715	=>	47081,
		4716	=>	47083,
		4717	=>	47086,
		4718	=>	47089,
		4719	=>	47092,
		4720	=>	47095,
		4721	=>	47097,
		4722	=>	47100,
		4723	=>	47103,
		4724	=>	47106,
		4725	=>	47109,
		4726	=>	47112,
		4727	=>	47114,
		4728	=>	47117,
		4729	=>	47120,
		4730	=>	47123,
		4731	=>	47126,
		4732	=>	47129,
		4733	=>	47131,
		4734	=>	47134,
		4735	=>	47137,
		4736	=>	47140,
		4737	=>	47143,
		4738	=>	47146,
		4739	=>	47148,
		4740	=>	47151,
		4741	=>	47154,
		4742	=>	47157,
		4743	=>	47160,
		4744	=>	47162,
		4745	=>	47165,
		4746	=>	47168,
		4747	=>	47171,
		4748	=>	47174,
		4749	=>	47177,
		4750	=>	47179,
		4751	=>	47182,
		4752	=>	47185,
		4753	=>	47188,
		4754	=>	47191,
		4755	=>	47193,
		4756	=>	47196,
		4757	=>	47199,
		4758	=>	47202,
		4759	=>	47205,
		4760	=>	47208,
		4761	=>	47210,
		4762	=>	47213,
		4763	=>	47216,
		4764	=>	47219,
		4765	=>	47222,
		4766	=>	47224,
		4767	=>	47227,
		4768	=>	47230,
		4769	=>	47233,
		4770	=>	47236,
		4771	=>	47239,
		4772	=>	47241,
		4773	=>	47244,
		4774	=>	47247,
		4775	=>	47250,
		4776	=>	47253,
		4777	=>	47255,
		4778	=>	47258,
		4779	=>	47261,
		4780	=>	47264,
		4781	=>	47267,
		4782	=>	47270,
		4783	=>	47272,
		4784	=>	47275,
		4785	=>	47278,
		4786	=>	47281,
		4787	=>	47284,
		4788	=>	47286,
		4789	=>	47289,
		4790	=>	47292,
		4791	=>	47295,
		4792	=>	47298,
		4793	=>	47301,
		4794	=>	47303,
		4795	=>	47306,
		4796	=>	47309,
		4797	=>	47312,
		4798	=>	47315,
		4799	=>	47317,
		4800	=>	47320,
		4801	=>	47323,
		4802	=>	47326,
		4803	=>	47329,
		4804	=>	47332,
		4805	=>	47334,
		4806	=>	47337,
		4807	=>	47340,
		4808	=>	47343,
		4809	=>	47346,
		4810	=>	47348,
		4811	=>	47351,
		4812	=>	47354,
		4813	=>	47357,
		4814	=>	47360,
		4815	=>	47362,
		4816	=>	47365,
		4817	=>	47368,
		4818	=>	47371,
		4819	=>	47374,
		4820	=>	47377,
		4821	=>	47379,
		4822	=>	47382,
		4823	=>	47385,
		4824	=>	47388,
		4825	=>	47391,
		4826	=>	47393,
		4827	=>	47396,
		4828	=>	47399,
		4829	=>	47402,
		4830	=>	47405,
		4831	=>	47407,
		4832	=>	47410,
		4833	=>	47413,
		4834	=>	47416,
		4835	=>	47419,
		4836	=>	47422,
		4837	=>	47424,
		4838	=>	47427,
		4839	=>	47430,
		4840	=>	47433,
		4841	=>	47436,
		4842	=>	47438,
		4843	=>	47441,
		4844	=>	47444,
		4845	=>	47447,
		4846	=>	47450,
		4847	=>	47452,
		4848	=>	47455,
		4849	=>	47458,
		4850	=>	47461,
		4851	=>	47464,
		4852	=>	47466,
		4853	=>	47469,
		4854	=>	47472,
		4855	=>	47475,
		4856	=>	47478,
		4857	=>	47480,
		4858	=>	47483,
		4859	=>	47486,
		4860	=>	47489,
		4861	=>	47492,
		4862	=>	47495,
		4863	=>	47497,
		4864	=>	47500,
		4865	=>	47503,
		4866	=>	47506,
		4867	=>	47509,
		4868	=>	47511,
		4869	=>	47514,
		4870	=>	47517,
		4871	=>	47520,
		4872	=>	47523,
		4873	=>	47525,
		4874	=>	47528,
		4875	=>	47531,
		4876	=>	47534,
		4877	=>	47537,
		4878	=>	47539,
		4879	=>	47542,
		4880	=>	47545,
		4881	=>	47548,
		4882	=>	47551,
		4883	=>	47553,
		4884	=>	47556,
		4885	=>	47559,
		4886	=>	47562,
		4887	=>	47565,
		4888	=>	47567,
		4889	=>	47570,
		4890	=>	47573,
		4891	=>	47576,
		4892	=>	47579,
		4893	=>	47581,
		4894	=>	47584,
		4895	=>	47587,
		4896	=>	47590,
		4897	=>	47593,
		4898	=>	47595,
		4899	=>	47598,
		4900	=>	47601,
		4901	=>	47604,
		4902	=>	47607,
		4903	=>	47609,
		4904	=>	47612,
		4905	=>	47615,
		4906	=>	47618,
		4907	=>	47621,
		4908	=>	47623,
		4909	=>	47626,
		4910	=>	47629,
		4911	=>	47632,
		4912	=>	47635,
		4913	=>	47637,
		4914	=>	47640,
		4915	=>	47643,
		4916	=>	47646,
		4917	=>	47649,
		4918	=>	47651,
		4919	=>	47654,
		4920	=>	47657,
		4921	=>	47660,
		4922	=>	47663,
		4923	=>	47665,
		4924	=>	47668,
		4925	=>	47671,
		4926	=>	47674,
		4927	=>	47677,
		4928	=>	47679,
		4929	=>	47682,
		4930	=>	47685,
		4931	=>	47688,
		4932	=>	47691,
		4933	=>	47693,
		4934	=>	47696,
		4935	=>	47699,
		4936	=>	47702,
		4937	=>	47705,
		4938	=>	47707,
		4939	=>	47710,
		4940	=>	47713,
		4941	=>	47716,
		4942	=>	47719,
		4943	=>	47721,
		4944	=>	47724,
		4945	=>	47727,
		4946	=>	47730,
		4947	=>	47733,
		4948	=>	47735,
		4949	=>	47738,
		4950	=>	47741,
		4951	=>	47744,
		4952	=>	47747,
		4953	=>	47749,
		4954	=>	47752,
		4955	=>	47755,
		4956	=>	47758,
		4957	=>	47761,
		4958	=>	47763,
		4959	=>	47766,
		4960	=>	47769,
		4961	=>	47772,
		4962	=>	47774,
		4963	=>	47777,
		4964	=>	47780,
		4965	=>	47783,
		4966	=>	47786,
		4967	=>	47788,
		4968	=>	47791,
		4969	=>	47794,
		4970	=>	47797,
		4971	=>	47800,
		4972	=>	47802,
		4973	=>	47805,
		4974	=>	47808,
		4975	=>	47811,
		4976	=>	47814,
		4977	=>	47816,
		4978	=>	47819,
		4979	=>	47822,
		4980	=>	47825,
		4981	=>	47828,
		4982	=>	47830,
		4983	=>	47833,
		4984	=>	47836,
		4985	=>	47839,
		4986	=>	47841,
		4987	=>	47844,
		4988	=>	47847,
		4989	=>	47850,
		4990	=>	47853,
		4991	=>	47855,
		4992	=>	47858,
		4993	=>	47861,
		4994	=>	47864,
		4995	=>	47867,
		4996	=>	47869,
		4997	=>	47872,
		4998	=>	47875,
		4999	=>	47878,
		5000	=>	47881,
		5001	=>	47883,
		5002	=>	47886,
		5003	=>	47889,
		5004	=>	47892,
		5005	=>	47894,
		5006	=>	47897,
		5007	=>	47900,
		5008	=>	47903,
		5009	=>	47906,
		5010	=>	47908,
		5011	=>	47911,
		5012	=>	47914,
		5013	=>	47917,
		5014	=>	47920,
		5015	=>	47922,
		5016	=>	47925,
		5017	=>	47928,
		5018	=>	47931,
		5019	=>	47933,
		5020	=>	47936,
		5021	=>	47939,
		5022	=>	47942,
		5023	=>	47945,
		5024	=>	47947,
		5025	=>	47950,
		5026	=>	47953,
		5027	=>	47956,
		5028	=>	47959,
		5029	=>	47961,
		5030	=>	47964,
		5031	=>	47967,
		5032	=>	47970,
		5033	=>	47972,
		5034	=>	47975,
		5035	=>	47978,
		5036	=>	47981,
		5037	=>	47984,
		5038	=>	47986,
		5039	=>	47989,
		5040	=>	47992,
		5041	=>	47995,
		5042	=>	47997,
		5043	=>	48000,
		5044	=>	48003,
		5045	=>	48006,
		5046	=>	48009,
		5047	=>	48011,
		5048	=>	48014,
		5049	=>	48017,
		5050	=>	48020,
		5051	=>	48022,
		5052	=>	48025,
		5053	=>	48028,
		5054	=>	48031,
		5055	=>	48034,
		5056	=>	48036,
		5057	=>	48039,
		5058	=>	48042,
		5059	=>	48045,
		5060	=>	48048,
		5061	=>	48050,
		5062	=>	48053,
		5063	=>	48056,
		5064	=>	48059,
		5065	=>	48061,
		5066	=>	48064,
		5067	=>	48067,
		5068	=>	48070,
		5069	=>	48073,
		5070	=>	48075,
		5071	=>	48078,
		5072	=>	48081,
		5073	=>	48084,
		5074	=>	48086,
		5075	=>	48089,
		5076	=>	48092,
		5077	=>	48095,
		5078	=>	48098,
		5079	=>	48100,
		5080	=>	48103,
		5081	=>	48106,
		5082	=>	48109,
		5083	=>	48111,
		5084	=>	48114,
		5085	=>	48117,
		5086	=>	48120,
		5087	=>	48122,
		5088	=>	48125,
		5089	=>	48128,
		5090	=>	48131,
		5091	=>	48134,
		5092	=>	48136,
		5093	=>	48139,
		5094	=>	48142,
		5095	=>	48145,
		5096	=>	48147,
		5097	=>	48150,
		5098	=>	48153,
		5099	=>	48156,
		5100	=>	48159,
		5101	=>	48161,
		5102	=>	48164,
		5103	=>	48167,
		5104	=>	48170,
		5105	=>	48172,
		5106	=>	48175,
		5107	=>	48178,
		5108	=>	48181,
		5109	=>	48184,
		5110	=>	48186,
		5111	=>	48189,
		5112	=>	48192,
		5113	=>	48195,
		5114	=>	48197,
		5115	=>	48200,
		5116	=>	48203,
		5117	=>	48206,
		5118	=>	48208,
		5119	=>	48211,
		5120	=>	48214,
		5121	=>	48217,
		5122	=>	48220,
		5123	=>	48222,
		5124	=>	48225,
		5125	=>	48228,
		5126	=>	48231,
		5127	=>	48233,
		5128	=>	48236,
		5129	=>	48239,
		5130	=>	48242,
		5131	=>	48244,
		5132	=>	48247,
		5133	=>	48250,
		5134	=>	48253,
		5135	=>	48256,
		5136	=>	48258,
		5137	=>	48261,
		5138	=>	48264,
		5139	=>	48267,
		5140	=>	48269,
		5141	=>	48272,
		5142	=>	48275,
		5143	=>	48278,
		5144	=>	48280,
		5145	=>	48283,
		5146	=>	48286,
		5147	=>	48289,
		5148	=>	48292,
		5149	=>	48294,
		5150	=>	48297,
		5151	=>	48300,
		5152	=>	48303,
		5153	=>	48305,
		5154	=>	48308,
		5155	=>	48311,
		5156	=>	48314,
		5157	=>	48316,
		5158	=>	48319,
		5159	=>	48322,
		5160	=>	48325,
		5161	=>	48327,
		5162	=>	48330,
		5163	=>	48333,
		5164	=>	48336,
		5165	=>	48339,
		5166	=>	48341,
		5167	=>	48344,
		5168	=>	48347,
		5169	=>	48350,
		5170	=>	48352,
		5171	=>	48355,
		5172	=>	48358,
		5173	=>	48361,
		5174	=>	48363,
		5175	=>	48366,
		5176	=>	48369,
		5177	=>	48372,
		5178	=>	48374,
		5179	=>	48377,
		5180	=>	48380,
		5181	=>	48383,
		5182	=>	48385,
		5183	=>	48388,
		5184	=>	48391,
		5185	=>	48394,
		5186	=>	48397,
		5187	=>	48399,
		5188	=>	48402,
		5189	=>	48405,
		5190	=>	48408,
		5191	=>	48410,
		5192	=>	48413,
		5193	=>	48416,
		5194	=>	48419,
		5195	=>	48421,
		5196	=>	48424,
		5197	=>	48427,
		5198	=>	48430,
		5199	=>	48432,
		5200	=>	48435,
		5201	=>	48438,
		5202	=>	48441,
		5203	=>	48443,
		5204	=>	48446,
		5205	=>	48449,
		5206	=>	48452,
		5207	=>	48454,
		5208	=>	48457,
		5209	=>	48460,
		5210	=>	48463,
		5211	=>	48466,
		5212	=>	48468,
		5213	=>	48471,
		5214	=>	48474,
		5215	=>	48477,
		5216	=>	48479,
		5217	=>	48482,
		5218	=>	48485,
		5219	=>	48488,
		5220	=>	48490,
		5221	=>	48493,
		5222	=>	48496,
		5223	=>	48499,
		5224	=>	48501,
		5225	=>	48504,
		5226	=>	48507,
		5227	=>	48510,
		5228	=>	48512,
		5229	=>	48515,
		5230	=>	48518,
		5231	=>	48521,
		5232	=>	48523,
		5233	=>	48526,
		5234	=>	48529,
		5235	=>	48532,
		5236	=>	48534,
		5237	=>	48537,
		5238	=>	48540,
		5239	=>	48543,
		5240	=>	48545,
		5241	=>	48548,
		5242	=>	48551,
		5243	=>	48554,
		5244	=>	48556,
		5245	=>	48559,
		5246	=>	48562,
		5247	=>	48565,
		5248	=>	48567,
		5249	=>	48570,
		5250	=>	48573,
		5251	=>	48576,
		5252	=>	48578,
		5253	=>	48581,
		5254	=>	48584,
		5255	=>	48587,
		5256	=>	48589,
		5257	=>	48592,
		5258	=>	48595,
		5259	=>	48598,
		5260	=>	48600,
		5261	=>	48603,
		5262	=>	48606,
		5263	=>	48609,
		5264	=>	48611,
		5265	=>	48614,
		5266	=>	48617,
		5267	=>	48620,
		5268	=>	48622,
		5269	=>	48625,
		5270	=>	48628,
		5271	=>	48631,
		5272	=>	48633,
		5273	=>	48636,
		5274	=>	48639,
		5275	=>	48642,
		5276	=>	48644,
		5277	=>	48647,
		5278	=>	48650,
		5279	=>	48653,
		5280	=>	48655,
		5281	=>	48658,
		5282	=>	48661,
		5283	=>	48664,
		5284	=>	48666,
		5285	=>	48669,
		5286	=>	48672,
		5287	=>	48675,
		5288	=>	48677,
		5289	=>	48680,
		5290	=>	48683,
		5291	=>	48686,
		5292	=>	48688,
		5293	=>	48691,
		5294	=>	48694,
		5295	=>	48697,
		5296	=>	48699,
		5297	=>	48702,
		5298	=>	48705,
		5299	=>	48708,
		5300	=>	48710,
		5301	=>	48713,
		5302	=>	48716,
		5303	=>	48719,
		5304	=>	48721,
		5305	=>	48724,
		5306	=>	48727,
		5307	=>	48730,
		5308	=>	48732,
		5309	=>	48735,
		5310	=>	48738,
		5311	=>	48741,
		5312	=>	48743,
		5313	=>	48746,
		5314	=>	48749,
		5315	=>	48752,
		5316	=>	48754,
		5317	=>	48757,
		5318	=>	48760,
		5319	=>	48762,
		5320	=>	48765,
		5321	=>	48768,
		5322	=>	48771,
		5323	=>	48773,
		5324	=>	48776,
		5325	=>	48779,
		5326	=>	48782,
		5327	=>	48784,
		5328	=>	48787,
		5329	=>	48790,
		5330	=>	48793,
		5331	=>	48795,
		5332	=>	48798,
		5333	=>	48801,
		5334	=>	48804,
		5335	=>	48806,
		5336	=>	48809,
		5337	=>	48812,
		5338	=>	48815,
		5339	=>	48817,
		5340	=>	48820,
		5341	=>	48823,
		5342	=>	48826,
		5343	=>	48828,
		5344	=>	48831,
		5345	=>	48834,
		5346	=>	48836,
		5347	=>	48839,
		5348	=>	48842,
		5349	=>	48845,
		5350	=>	48847,
		5351	=>	48850,
		5352	=>	48853,
		5353	=>	48856,
		5354	=>	48858,
		5355	=>	48861,
		5356	=>	48864,
		5357	=>	48867,
		5358	=>	48869,
		5359	=>	48872,
		5360	=>	48875,
		5361	=>	48878,
		5362	=>	48880,
		5363	=>	48883,
		5364	=>	48886,
		5365	=>	48888,
		5366	=>	48891,
		5367	=>	48894,
		5368	=>	48897,
		5369	=>	48899,
		5370	=>	48902,
		5371	=>	48905,
		5372	=>	48908,
		5373	=>	48910,
		5374	=>	48913,
		5375	=>	48916,
		5376	=>	48919,
		5377	=>	48921,
		5378	=>	48924,
		5379	=>	48927,
		5380	=>	48929,
		5381	=>	48932,
		5382	=>	48935,
		5383	=>	48938,
		5384	=>	48940,
		5385	=>	48943,
		5386	=>	48946,
		5387	=>	48949,
		5388	=>	48951,
		5389	=>	48954,
		5390	=>	48957,
		5391	=>	48960,
		5392	=>	48962,
		5393	=>	48965,
		5394	=>	48968,
		5395	=>	48970,
		5396	=>	48973,
		5397	=>	48976,
		5398	=>	48979,
		5399	=>	48981,
		5400	=>	48984,
		5401	=>	48987,
		5402	=>	48990,
		5403	=>	48992,
		5404	=>	48995,
		5405	=>	48998,
		5406	=>	49000,
		5407	=>	49003,
		5408	=>	49006,
		5409	=>	49009,
		5410	=>	49011,
		5411	=>	49014,
		5412	=>	49017,
		5413	=>	49020,
		5414	=>	49022,
		5415	=>	49025,
		5416	=>	49028,
		5417	=>	49030,
		5418	=>	49033,
		5419	=>	49036,
		5420	=>	49039,
		5421	=>	49041,
		5422	=>	49044,
		5423	=>	49047,
		5424	=>	49050,
		5425	=>	49052,
		5426	=>	49055,
		5427	=>	49058,
		5428	=>	49060,
		5429	=>	49063,
		5430	=>	49066,
		5431	=>	49069,
		5432	=>	49071,
		5433	=>	49074,
		5434	=>	49077,
		5435	=>	49080,
		5436	=>	49082,
		5437	=>	49085,
		5438	=>	49088,
		5439	=>	49090,
		5440	=>	49093,
		5441	=>	49096,
		5442	=>	49099,
		5443	=>	49101,
		5444	=>	49104,
		5445	=>	49107,
		5446	=>	49110,
		5447	=>	49112,
		5448	=>	49115,
		5449	=>	49118,
		5450	=>	49120,
		5451	=>	49123,
		5452	=>	49126,
		5453	=>	49129,
		5454	=>	49131,
		5455	=>	49134,
		5456	=>	49137,
		5457	=>	49139,
		5458	=>	49142,
		5459	=>	49145,
		5460	=>	49148,
		5461	=>	49150,
		5462	=>	49153,
		5463	=>	49156,
		5464	=>	49159,
		5465	=>	49161,
		5466	=>	49164,
		5467	=>	49167,
		5468	=>	49169,
		5469	=>	49172,
		5470	=>	49175,
		5471	=>	49178,
		5472	=>	49180,
		5473	=>	49183,
		5474	=>	49186,
		5475	=>	49188,
		5476	=>	49191,
		5477	=>	49194,
		5478	=>	49197,
		5479	=>	49199,
		5480	=>	49202,
		5481	=>	49205,
		5482	=>	49207,
		5483	=>	49210,
		5484	=>	49213,
		5485	=>	49216,
		5486	=>	49218,
		5487	=>	49221,
		5488	=>	49224,
		5489	=>	49226,
		5490	=>	49229,
		5491	=>	49232,
		5492	=>	49235,
		5493	=>	49237,
		5494	=>	49240,
		5495	=>	49243,
		5496	=>	49245,
		5497	=>	49248,
		5498	=>	49251,
		5499	=>	49254,
		5500	=>	49256,
		5501	=>	49259,
		5502	=>	49262,
		5503	=>	49264,
		5504	=>	49267,
		5505	=>	49270,
		5506	=>	49273,
		5507	=>	49275,
		5508	=>	49278,
		5509	=>	49281,
		5510	=>	49283,
		5511	=>	49286,
		5512	=>	49289,
		5513	=>	49292,
		5514	=>	49294,
		5515	=>	49297,
		5516	=>	49300,
		5517	=>	49302,
		5518	=>	49305,
		5519	=>	49308,
		5520	=>	49311,
		5521	=>	49313,
		5522	=>	49316,
		5523	=>	49319,
		5524	=>	49321,
		5525	=>	49324,
		5526	=>	49327,
		5527	=>	49330,
		5528	=>	49332,
		5529	=>	49335,
		5530	=>	49338,
		5531	=>	49340,
		5532	=>	49343,
		5533	=>	49346,
		5534	=>	49349,
		5535	=>	49351,
		5536	=>	49354,
		5537	=>	49357,
		5538	=>	49359,
		5539	=>	49362,
		5540	=>	49365,
		5541	=>	49368,
		5542	=>	49370,
		5543	=>	49373,
		5544	=>	49376,
		5545	=>	49378,
		5546	=>	49381,
		5547	=>	49384,
		5548	=>	49386,
		5549	=>	49389,
		5550	=>	49392,
		5551	=>	49395,
		5552	=>	49397,
		5553	=>	49400,
		5554	=>	49403,
		5555	=>	49405,
		5556	=>	49408,
		5557	=>	49411,
		5558	=>	49414,
		5559	=>	49416,
		5560	=>	49419,
		5561	=>	49422,
		5562	=>	49424,
		5563	=>	49427,
		5564	=>	49430,
		5565	=>	49432,
		5566	=>	49435,
		5567	=>	49438,
		5568	=>	49441,
		5569	=>	49443,
		5570	=>	49446,
		5571	=>	49449,
		5572	=>	49451,
		5573	=>	49454,
		5574	=>	49457,
		5575	=>	49460,
		5576	=>	49462,
		5577	=>	49465,
		5578	=>	49468,
		5579	=>	49470,
		5580	=>	49473,
		5581	=>	49476,
		5582	=>	49478,
		5583	=>	49481,
		5584	=>	49484,
		5585	=>	49487,
		5586	=>	49489,
		5587	=>	49492,
		5588	=>	49495,
		5589	=>	49497,
		5590	=>	49500,
		5591	=>	49503,
		5592	=>	49505,
		5593	=>	49508,
		5594	=>	49511,
		5595	=>	49514,
		5596	=>	49516,
		5597	=>	49519,
		5598	=>	49522,
		5599	=>	49524,
		5600	=>	49527,
		5601	=>	49530,
		5602	=>	49532,
		5603	=>	49535,
		5604	=>	49538,
		5605	=>	49541,
		5606	=>	49543,
		5607	=>	49546,
		5608	=>	49549,
		5609	=>	49551,
		5610	=>	49554,
		5611	=>	49557,
		5612	=>	49559,
		5613	=>	49562,
		5614	=>	49565,
		5615	=>	49568,
		5616	=>	49570,
		5617	=>	49573,
		5618	=>	49576,
		5619	=>	49578,
		5620	=>	49581,
		5621	=>	49584,
		5622	=>	49586,
		5623	=>	49589,
		5624	=>	49592,
		5625	=>	49594,
		5626	=>	49597,
		5627	=>	49600,
		5628	=>	49603,
		5629	=>	49605,
		5630	=>	49608,
		5631	=>	49611,
		5632	=>	49613,
		5633	=>	49616,
		5634	=>	49619,
		5635	=>	49621,
		5636	=>	49624,
		5637	=>	49627,
		5638	=>	49630,
		5639	=>	49632,
		5640	=>	49635,
		5641	=>	49638,
		5642	=>	49640,
		5643	=>	49643,
		5644	=>	49646,
		5645	=>	49648,
		5646	=>	49651,
		5647	=>	49654,
		5648	=>	49656,
		5649	=>	49659,
		5650	=>	49662,
		5651	=>	49665,
		5652	=>	49667,
		5653	=>	49670,
		5654	=>	49673,
		5655	=>	49675,
		5656	=>	49678,
		5657	=>	49681,
		5658	=>	49683,
		5659	=>	49686,
		5660	=>	49689,
		5661	=>	49691,
		5662	=>	49694,
		5663	=>	49697,
		5664	=>	49700,
		5665	=>	49702,
		5666	=>	49705,
		5667	=>	49708,
		5668	=>	49710,
		5669	=>	49713,
		5670	=>	49716,
		5671	=>	49718,
		5672	=>	49721,
		5673	=>	49724,
		5674	=>	49726,
		5675	=>	49729,
		5676	=>	49732,
		5677	=>	49734,
		5678	=>	49737,
		5679	=>	49740,
		5680	=>	49743,
		5681	=>	49745,
		5682	=>	49748,
		5683	=>	49751,
		5684	=>	49753,
		5685	=>	49756,
		5686	=>	49759,
		5687	=>	49761,
		5688	=>	49764,
		5689	=>	49767,
		5690	=>	49769,
		5691	=>	49772,
		5692	=>	49775,
		5693	=>	49777,
		5694	=>	49780,
		5695	=>	49783,
		5696	=>	49785,
		5697	=>	49788,
		5698	=>	49791,
		5699	=>	49794,
		5700	=>	49796,
		5701	=>	49799,
		5702	=>	49802,
		5703	=>	49804,
		5704	=>	49807,
		5705	=>	49810,
		5706	=>	49812,
		5707	=>	49815,
		5708	=>	49818,
		5709	=>	49820,
		5710	=>	49823,
		5711	=>	49826,
		5712	=>	49828,
		5713	=>	49831,
		5714	=>	49834,
		5715	=>	49836,
		5716	=>	49839,
		5717	=>	49842,
		5718	=>	49845,
		5719	=>	49847,
		5720	=>	49850,
		5721	=>	49853,
		5722	=>	49855,
		5723	=>	49858,
		5724	=>	49861,
		5725	=>	49863,
		5726	=>	49866,
		5727	=>	49869,
		5728	=>	49871,
		5729	=>	49874,
		5730	=>	49877,
		5731	=>	49879,
		5732	=>	49882,
		5733	=>	49885,
		5734	=>	49887,
		5735	=>	49890,
		5736	=>	49893,
		5737	=>	49895,
		5738	=>	49898,
		5739	=>	49901,
		5740	=>	49903,
		5741	=>	49906,
		5742	=>	49909,
		5743	=>	49912,
		5744	=>	49914,
		5745	=>	49917,
		5746	=>	49920,
		5747	=>	49922,
		5748	=>	49925,
		5749	=>	49928,
		5750	=>	49930,
		5751	=>	49933,
		5752	=>	49936,
		5753	=>	49938,
		5754	=>	49941,
		5755	=>	49944,
		5756	=>	49946,
		5757	=>	49949,
		5758	=>	49952,
		5759	=>	49954,
		5760	=>	49957,
		5761	=>	49960,
		5762	=>	49962,
		5763	=>	49965,
		5764	=>	49968,
		5765	=>	49970,
		5766	=>	49973,
		5767	=>	49976,
		5768	=>	49978,
		5769	=>	49981,
		5770	=>	49984,
		5771	=>	49986,
		5772	=>	49989,
		5773	=>	49992,
		5774	=>	49994,
		5775	=>	49997,
		5776	=>	50000,
		5777	=>	50002,
		5778	=>	50005,
		5779	=>	50008,
		5780	=>	50010,
		5781	=>	50013,
		5782	=>	50016,
		5783	=>	50018,
		5784	=>	50021,
		5785	=>	50024,
		5786	=>	50026,
		5787	=>	50029,
		5788	=>	50032,
		5789	=>	50034,
		5790	=>	50037,
		5791	=>	50040,
		5792	=>	50042,
		5793	=>	50045,
		5794	=>	50048,
		5795	=>	50051,
		5796	=>	50053,
		5797	=>	50056,
		5798	=>	50059,
		5799	=>	50061,
		5800	=>	50064,
		5801	=>	50067,
		5802	=>	50069,
		5803	=>	50072,
		5804	=>	50075,
		5805	=>	50077,
		5806	=>	50080,
		5807	=>	50083,
		5808	=>	50085,
		5809	=>	50088,
		5810	=>	50091,
		5811	=>	50093,
		5812	=>	50096,
		5813	=>	50099,
		5814	=>	50101,
		5815	=>	50104,
		5816	=>	50107,
		5817	=>	50109,
		5818	=>	50112,
		5819	=>	50115,
		5820	=>	50117,
		5821	=>	50120,
		5822	=>	50123,
		5823	=>	50125,
		5824	=>	50128,
		5825	=>	50131,
		5826	=>	50133,
		5827	=>	50136,
		5828	=>	50138,
		5829	=>	50141,
		5830	=>	50144,
		5831	=>	50146,
		5832	=>	50149,
		5833	=>	50152,
		5834	=>	50154,
		5835	=>	50157,
		5836	=>	50160,
		5837	=>	50162,
		5838	=>	50165,
		5839	=>	50168,
		5840	=>	50170,
		5841	=>	50173,
		5842	=>	50176,
		5843	=>	50178,
		5844	=>	50181,
		5845	=>	50184,
		5846	=>	50186,
		5847	=>	50189,
		5848	=>	50192,
		5849	=>	50194,
		5850	=>	50197,
		5851	=>	50200,
		5852	=>	50202,
		5853	=>	50205,
		5854	=>	50208,
		5855	=>	50210,
		5856	=>	50213,
		5857	=>	50216,
		5858	=>	50218,
		5859	=>	50221,
		5860	=>	50224,
		5861	=>	50226,
		5862	=>	50229,
		5863	=>	50232,
		5864	=>	50234,
		5865	=>	50237,
		5866	=>	50240,
		5867	=>	50242,
		5868	=>	50245,
		5869	=>	50248,
		5870	=>	50250,
		5871	=>	50253,
		5872	=>	50256,
		5873	=>	50258,
		5874	=>	50261,
		5875	=>	50264,
		5876	=>	50266,
		5877	=>	50269,
		5878	=>	50271,
		5879	=>	50274,
		5880	=>	50277,
		5881	=>	50279,
		5882	=>	50282,
		5883	=>	50285,
		5884	=>	50287,
		5885	=>	50290,
		5886	=>	50293,
		5887	=>	50295,
		5888	=>	50298,
		5889	=>	50301,
		5890	=>	50303,
		5891	=>	50306,
		5892	=>	50309,
		5893	=>	50311,
		5894	=>	50314,
		5895	=>	50317,
		5896	=>	50319,
		5897	=>	50322,
		5898	=>	50325,
		5899	=>	50327,
		5900	=>	50330,
		5901	=>	50333,
		5902	=>	50335,
		5903	=>	50338,
		5904	=>	50340,
		5905	=>	50343,
		5906	=>	50346,
		5907	=>	50348,
		5908	=>	50351,
		5909	=>	50354,
		5910	=>	50356,
		5911	=>	50359,
		5912	=>	50362,
		5913	=>	50364,
		5914	=>	50367,
		5915	=>	50370,
		5916	=>	50372,
		5917	=>	50375,
		5918	=>	50378,
		5919	=>	50380,
		5920	=>	50383,
		5921	=>	50386,
		5922	=>	50388,
		5923	=>	50391,
		5924	=>	50393,
		5925	=>	50396,
		5926	=>	50399,
		5927	=>	50401,
		5928	=>	50404,
		5929	=>	50407,
		5930	=>	50409,
		5931	=>	50412,
		5932	=>	50415,
		5933	=>	50417,
		5934	=>	50420,
		5935	=>	50423,
		5936	=>	50425,
		5937	=>	50428,
		5938	=>	50431,
		5939	=>	50433,
		5940	=>	50436,
		5941	=>	50438,
		5942	=>	50441,
		5943	=>	50444,
		5944	=>	50446,
		5945	=>	50449,
		5946	=>	50452,
		5947	=>	50454,
		5948	=>	50457,
		5949	=>	50460,
		5950	=>	50462,
		5951	=>	50465,
		5952	=>	50468,
		5953	=>	50470,
		5954	=>	50473,
		5955	=>	50475,
		5956	=>	50478,
		5957	=>	50481,
		5958	=>	50483,
		5959	=>	50486,
		5960	=>	50489,
		5961	=>	50491,
		5962	=>	50494,
		5963	=>	50497,
		5964	=>	50499,
		5965	=>	50502,
		5966	=>	50505,
		5967	=>	50507,
		5968	=>	50510,
		5969	=>	50512,
		5970	=>	50515,
		5971	=>	50518,
		5972	=>	50520,
		5973	=>	50523,
		5974	=>	50526,
		5975	=>	50528,
		5976	=>	50531,
		5977	=>	50534,
		5978	=>	50536,
		5979	=>	50539,
		5980	=>	50542,
		5981	=>	50544,
		5982	=>	50547,
		5983	=>	50549,
		5984	=>	50552,
		5985	=>	50555,
		5986	=>	50557,
		5987	=>	50560,
		5988	=>	50563,
		5989	=>	50565,
		5990	=>	50568,
		5991	=>	50571,
		5992	=>	50573,
		5993	=>	50576,
		5994	=>	50578,
		5995	=>	50581,
		5996	=>	50584,
		5997	=>	50586,
		5998	=>	50589,
		5999	=>	50592,
		6000	=>	50594,
		6001	=>	50597,
		6002	=>	50600,
		6003	=>	50602,
		6004	=>	50605,
		6005	=>	50607,
		6006	=>	50610,
		6007	=>	50613,
		6008	=>	50615,
		6009	=>	50618,
		6010	=>	50621,
		6011	=>	50623,
		6012	=>	50626,
		6013	=>	50629,
		6014	=>	50631,
		6015	=>	50634,
		6016	=>	50636,
		6017	=>	50639,
		6018	=>	50642,
		6019	=>	50644,
		6020	=>	50647,
		6021	=>	50650,
		6022	=>	50652,
		6023	=>	50655,
		6024	=>	50657,
		6025	=>	50660,
		6026	=>	50663,
		6027	=>	50665,
		6028	=>	50668,
		6029	=>	50671,
		6030	=>	50673,
		6031	=>	50676,
		6032	=>	50679,
		6033	=>	50681,
		6034	=>	50684,
		6035	=>	50686,
		6036	=>	50689,
		6037	=>	50692,
		6038	=>	50694,
		6039	=>	50697,
		6040	=>	50700,
		6041	=>	50702,
		6042	=>	50705,
		6043	=>	50707,
		6044	=>	50710,
		6045	=>	50713,
		6046	=>	50715,
		6047	=>	50718,
		6048	=>	50721,
		6049	=>	50723,
		6050	=>	50726,
		6051	=>	50729,
		6052	=>	50731,
		6053	=>	50734,
		6054	=>	50736,
		6055	=>	50739,
		6056	=>	50742,
		6057	=>	50744,
		6058	=>	50747,
		6059	=>	50750,
		6060	=>	50752,
		6061	=>	50755,
		6062	=>	50757,
		6063	=>	50760,
		6064	=>	50763,
		6065	=>	50765,
		6066	=>	50768,
		6067	=>	50771,
		6068	=>	50773,
		6069	=>	50776,
		6070	=>	50778,
		6071	=>	50781,
		6072	=>	50784,
		6073	=>	50786,
		6074	=>	50789,
		6075	=>	50792,
		6076	=>	50794,
		6077	=>	50797,
		6078	=>	50799,
		6079	=>	50802,
		6080	=>	50805,
		6081	=>	50807,
		6082	=>	50810,
		6083	=>	50812,
		6084	=>	50815,
		6085	=>	50818,
		6086	=>	50820,
		6087	=>	50823,
		6088	=>	50826,
		6089	=>	50828,
		6090	=>	50831,
		6091	=>	50833,
		6092	=>	50836,
		6093	=>	50839,
		6094	=>	50841,
		6095	=>	50844,
		6096	=>	50847,
		6097	=>	50849,
		6098	=>	50852,
		6099	=>	50854,
		6100	=>	50857,
		6101	=>	50860,
		6102	=>	50862,
		6103	=>	50865,
		6104	=>	50868,
		6105	=>	50870,
		6106	=>	50873,
		6107	=>	50875,
		6108	=>	50878,
		6109	=>	50881,
		6110	=>	50883,
		6111	=>	50886,
		6112	=>	50888,
		6113	=>	50891,
		6114	=>	50894,
		6115	=>	50896,
		6116	=>	50899,
		6117	=>	50902,
		6118	=>	50904,
		6119	=>	50907,
		6120	=>	50909,
		6121	=>	50912,
		6122	=>	50915,
		6123	=>	50917,
		6124	=>	50920,
		6125	=>	50922,
		6126	=>	50925,
		6127	=>	50928,
		6128	=>	50930,
		6129	=>	50933,
		6130	=>	50936,
		6131	=>	50938,
		6132	=>	50941,
		6133	=>	50943,
		6134	=>	50946,
		6135	=>	50949,
		6136	=>	50951,
		6137	=>	50954,
		6138	=>	50956,
		6139	=>	50959,
		6140	=>	50962,
		6141	=>	50964,
		6142	=>	50967,
		6143	=>	50970,
		6144	=>	50972,
		6145	=>	50975,
		6146	=>	50977,
		6147	=>	50980,
		6148	=>	50983,
		6149	=>	50985,
		6150	=>	50988,
		6151	=>	50990,
		6152	=>	50993,
		6153	=>	50996,
		6154	=>	50998,
		6155	=>	51001,
		6156	=>	51003,
		6157	=>	51006,
		6158	=>	51009,
		6159	=>	51011,
		6160	=>	51014,
		6161	=>	51017,
		6162	=>	51019,
		6163	=>	51022,
		6164	=>	51024,
		6165	=>	51027,
		6166	=>	51030,
		6167	=>	51032,
		6168	=>	51035,
		6169	=>	51037,
		6170	=>	51040,
		6171	=>	51043,
		6172	=>	51045,
		6173	=>	51048,
		6174	=>	51050,
		6175	=>	51053,
		6176	=>	51056,
		6177	=>	51058,
		6178	=>	51061,
		6179	=>	51063,
		6180	=>	51066,
		6181	=>	51069,
		6182	=>	51071,
		6183	=>	51074,
		6184	=>	51076,
		6185	=>	51079,
		6186	=>	51082,
		6187	=>	51084,
		6188	=>	51087,
		6189	=>	51090,
		6190	=>	51092,
		6191	=>	51095,
		6192	=>	51097,
		6193	=>	51100,
		6194	=>	51103,
		6195	=>	51105,
		6196	=>	51108,
		6197	=>	51110,
		6198	=>	51113,
		6199	=>	51116,
		6200	=>	51118,
		6201	=>	51121,
		6202	=>	51123,
		6203	=>	51126,
		6204	=>	51129,
		6205	=>	51131,
		6206	=>	51134,
		6207	=>	51136,
		6208	=>	51139,
		6209	=>	51142,
		6210	=>	51144,
		6211	=>	51147,
		6212	=>	51149,
		6213	=>	51152,
		6214	=>	51155,
		6215	=>	51157,
		6216	=>	51160,
		6217	=>	51162,
		6218	=>	51165,
		6219	=>	51168,
		6220	=>	51170,
		6221	=>	51173,
		6222	=>	51175,
		6223	=>	51178,
		6224	=>	51181,
		6225	=>	51183,
		6226	=>	51186,
		6227	=>	51188,
		6228	=>	51191,
		6229	=>	51194,
		6230	=>	51196,
		6231	=>	51199,
		6232	=>	51201,
		6233	=>	51204,
		6234	=>	51207,
		6235	=>	51209,
		6236	=>	51212,
		6237	=>	51214,
		6238	=>	51217,
		6239	=>	51220,
		6240	=>	51222,
		6241	=>	51225,
		6242	=>	51227,
		6243	=>	51230,
		6244	=>	51233,
		6245	=>	51235,
		6246	=>	51238,
		6247	=>	51240,
		6248	=>	51243,
		6249	=>	51245,
		6250	=>	51248,
		6251	=>	51251,
		6252	=>	51253,
		6253	=>	51256,
		6254	=>	51258,
		6255	=>	51261,
		6256	=>	51264,
		6257	=>	51266,
		6258	=>	51269,
		6259	=>	51271,
		6260	=>	51274,
		6261	=>	51277,
		6262	=>	51279,
		6263	=>	51282,
		6264	=>	51284,
		6265	=>	51287,
		6266	=>	51290,
		6267	=>	51292,
		6268	=>	51295,
		6269	=>	51297,
		6270	=>	51300,
		6271	=>	51303,
		6272	=>	51305,
		6273	=>	51308,
		6274	=>	51310,
		6275	=>	51313,
		6276	=>	51315,
		6277	=>	51318,
		6278	=>	51321,
		6279	=>	51323,
		6280	=>	51326,
		6281	=>	51328,
		6282	=>	51331,
		6283	=>	51334,
		6284	=>	51336,
		6285	=>	51339,
		6286	=>	51341,
		6287	=>	51344,
		6288	=>	51347,
		6289	=>	51349,
		6290	=>	51352,
		6291	=>	51354,
		6292	=>	51357,
		6293	=>	51359,
		6294	=>	51362,
		6295	=>	51365,
		6296	=>	51367,
		6297	=>	51370,
		6298	=>	51372,
		6299	=>	51375,
		6300	=>	51378,
		6301	=>	51380,
		6302	=>	51383,
		6303	=>	51385,
		6304	=>	51388,
		6305	=>	51391,
		6306	=>	51393,
		6307	=>	51396,
		6308	=>	51398,
		6309	=>	51401,
		6310	=>	51403,
		6311	=>	51406,
		6312	=>	51409,
		6313	=>	51411,
		6314	=>	51414,
		6315	=>	51416,
		6316	=>	51419,
		6317	=>	51422,
		6318	=>	51424,
		6319	=>	51427,
		6320	=>	51429,
		6321	=>	51432,
		6322	=>	51434,
		6323	=>	51437,
		6324	=>	51440,
		6325	=>	51442,
		6326	=>	51445,
		6327	=>	51447,
		6328	=>	51450,
		6329	=>	51452,
		6330	=>	51455,
		6331	=>	51458,
		6332	=>	51460,
		6333	=>	51463,
		6334	=>	51465,
		6335	=>	51468,
		6336	=>	51471,
		6337	=>	51473,
		6338	=>	51476,
		6339	=>	51478,
		6340	=>	51481,
		6341	=>	51483,
		6342	=>	51486,
		6343	=>	51489,
		6344	=>	51491,
		6345	=>	51494,
		6346	=>	51496,
		6347	=>	51499,
		6348	=>	51502,
		6349	=>	51504,
		6350	=>	51507,
		6351	=>	51509,
		6352	=>	51512,
		6353	=>	51514,
		6354	=>	51517,
		6355	=>	51520,
		6356	=>	51522,
		6357	=>	51525,
		6358	=>	51527,
		6359	=>	51530,
		6360	=>	51532,
		6361	=>	51535,
		6362	=>	51538,
		6363	=>	51540,
		6364	=>	51543,
		6365	=>	51545,
		6366	=>	51548,
		6367	=>	51550,
		6368	=>	51553,
		6369	=>	51556,
		6370	=>	51558,
		6371	=>	51561,
		6372	=>	51563,
		6373	=>	51566,
		6374	=>	51568,
		6375	=>	51571,
		6376	=>	51574,
		6377	=>	51576,
		6378	=>	51579,
		6379	=>	51581,
		6380	=>	51584,
		6381	=>	51586,
		6382	=>	51589,
		6383	=>	51592,
		6384	=>	51594,
		6385	=>	51597,
		6386	=>	51599,
		6387	=>	51602,
		6388	=>	51604,
		6389	=>	51607,
		6390	=>	51610,
		6391	=>	51612,
		6392	=>	51615,
		6393	=>	51617,
		6394	=>	51620,
		6395	=>	51622,
		6396	=>	51625,
		6397	=>	51628,
		6398	=>	51630,
		6399	=>	51633,
		6400	=>	51635,
		6401	=>	51638,
		6402	=>	51640,
		6403	=>	51643,
		6404	=>	51646,
		6405	=>	51648,
		6406	=>	51651,
		6407	=>	51653,
		6408	=>	51656,
		6409	=>	51658,
		6410	=>	51661,
		6411	=>	51664,
		6412	=>	51666,
		6413	=>	51669,
		6414	=>	51671,
		6415	=>	51674,
		6416	=>	51676,
		6417	=>	51679,
		6418	=>	51681,
		6419	=>	51684,
		6420	=>	51687,
		6421	=>	51689,
		6422	=>	51692,
		6423	=>	51694,
		6424	=>	51697,
		6425	=>	51699,
		6426	=>	51702,
		6427	=>	51705,
		6428	=>	51707,
		6429	=>	51710,
		6430	=>	51712,
		6431	=>	51715,
		6432	=>	51717,
		6433	=>	51720,
		6434	=>	51723,
		6435	=>	51725,
		6436	=>	51728,
		6437	=>	51730,
		6438	=>	51733,
		6439	=>	51735,
		6440	=>	51738,
		6441	=>	51740,
		6442	=>	51743,
		6443	=>	51746,
		6444	=>	51748,
		6445	=>	51751,
		6446	=>	51753,
		6447	=>	51756,
		6448	=>	51758,
		6449	=>	51761,
		6450	=>	51764,
		6451	=>	51766,
		6452	=>	51769,
		6453	=>	51771,
		6454	=>	51774,
		6455	=>	51776,
		6456	=>	51779,
		6457	=>	51781,
		6458	=>	51784,
		6459	=>	51787,
		6460	=>	51789,
		6461	=>	51792,
		6462	=>	51794,
		6463	=>	51797,
		6464	=>	51799,
		6465	=>	51802,
		6466	=>	51804,
		6467	=>	51807,
		6468	=>	51810,
		6469	=>	51812,
		6470	=>	51815,
		6471	=>	51817,
		6472	=>	51820,
		6473	=>	51822,
		6474	=>	51825,
		6475	=>	51827,
		6476	=>	51830,
		6477	=>	51833,
		6478	=>	51835,
		6479	=>	51838,
		6480	=>	51840,
		6481	=>	51843,
		6482	=>	51845,
		6483	=>	51848,
		6484	=>	51850,
		6485	=>	51853,
		6486	=>	51856,
		6487	=>	51858,
		6488	=>	51861,
		6489	=>	51863,
		6490	=>	51866,
		6491	=>	51868,
		6492	=>	51871,
		6493	=>	51873,
		6494	=>	51876,
		6495	=>	51879,
		6496	=>	51881,
		6497	=>	51884,
		6498	=>	51886,
		6499	=>	51889,
		6500	=>	51891,
		6501	=>	51894,
		6502	=>	51896,
		6503	=>	51899,
		6504	=>	51901,
		6505	=>	51904,
		6506	=>	51907,
		6507	=>	51909,
		6508	=>	51912,
		6509	=>	51914,
		6510	=>	51917,
		6511	=>	51919,
		6512	=>	51922,
		6513	=>	51924,
		6514	=>	51927,
		6515	=>	51930,
		6516	=>	51932,
		6517	=>	51935,
		6518	=>	51937,
		6519	=>	51940,
		6520	=>	51942,
		6521	=>	51945,
		6522	=>	51947,
		6523	=>	51950,
		6524	=>	51952,
		6525	=>	51955,
		6526	=>	51958,
		6527	=>	51960,
		6528	=>	51963,
		6529	=>	51965,
		6530	=>	51968,
		6531	=>	51970,
		6532	=>	51973,
		6533	=>	51975,
		6534	=>	51978,
		6535	=>	51980,
		6536	=>	51983,
		6537	=>	51986,
		6538	=>	51988,
		6539	=>	51991,
		6540	=>	51993,
		6541	=>	51996,
		6542	=>	51998,
		6543	=>	52001,
		6544	=>	52003,
		6545	=>	52006,
		6546	=>	52008,
		6547	=>	52011,
		6548	=>	52014,
		6549	=>	52016,
		6550	=>	52019,
		6551	=>	52021,
		6552	=>	52024,
		6553	=>	52026,
		6554	=>	52029,
		6555	=>	52031,
		6556	=>	52034,
		6557	=>	52036,
		6558	=>	52039,
		6559	=>	52041,
		6560	=>	52044,
		6561	=>	52047,
		6562	=>	52049,
		6563	=>	52052,
		6564	=>	52054,
		6565	=>	52057,
		6566	=>	52059,
		6567	=>	52062,
		6568	=>	52064,
		6569	=>	52067,
		6570	=>	52069,
		6571	=>	52072,
		6572	=>	52074,
		6573	=>	52077,
		6574	=>	52080,
		6575	=>	52082,
		6576	=>	52085,
		6577	=>	52087,
		6578	=>	52090,
		6579	=>	52092,
		6580	=>	52095,
		6581	=>	52097,
		6582	=>	52100,
		6583	=>	52102,
		6584	=>	52105,
		6585	=>	52107,
		6586	=>	52110,
		6587	=>	52113,
		6588	=>	52115,
		6589	=>	52118,
		6590	=>	52120,
		6591	=>	52123,
		6592	=>	52125,
		6593	=>	52128,
		6594	=>	52130,
		6595	=>	52133,
		6596	=>	52135,
		6597	=>	52138,
		6598	=>	52140,
		6599	=>	52143,
		6600	=>	52145,
		6601	=>	52148,
		6602	=>	52151,
		6603	=>	52153,
		6604	=>	52156,
		6605	=>	52158,
		6606	=>	52161,
		6607	=>	52163,
		6608	=>	52166,
		6609	=>	52168,
		6610	=>	52171,
		6611	=>	52173,
		6612	=>	52176,
		6613	=>	52178,
		6614	=>	52181,
		6615	=>	52183,
		6616	=>	52186,
		6617	=>	52189,
		6618	=>	52191,
		6619	=>	52194,
		6620	=>	52196,
		6621	=>	52199,
		6622	=>	52201,
		6623	=>	52204,
		6624	=>	52206,
		6625	=>	52209,
		6626	=>	52211,
		6627	=>	52214,
		6628	=>	52216,
		6629	=>	52219,
		6630	=>	52221,
		6631	=>	52224,
		6632	=>	52226,
		6633	=>	52229,
		6634	=>	52232,
		6635	=>	52234,
		6636	=>	52237,
		6637	=>	52239,
		6638	=>	52242,
		6639	=>	52244,
		6640	=>	52247,
		6641	=>	52249,
		6642	=>	52252,
		6643	=>	52254,
		6644	=>	52257,
		6645	=>	52259,
		6646	=>	52262,
		6647	=>	52264,
		6648	=>	52267,
		6649	=>	52269,
		6650	=>	52272,
		6651	=>	52274,
		6652	=>	52277,
		6653	=>	52280,
		6654	=>	52282,
		6655	=>	52285,
		6656	=>	52287,
		6657	=>	52290,
		6658	=>	52292,
		6659	=>	52295,
		6660	=>	52297,
		6661	=>	52300,
		6662	=>	52302,
		6663	=>	52305,
		6664	=>	52307,
		6665	=>	52310,
		6666	=>	52312,
		6667	=>	52315,
		6668	=>	52317,
		6669	=>	52320,
		6670	=>	52322,
		6671	=>	52325,
		6672	=>	52327,
		6673	=>	52330,
		6674	=>	52332,
		6675	=>	52335,
		6676	=>	52338,
		6677	=>	52340,
		6678	=>	52343,
		6679	=>	52345,
		6680	=>	52348,
		6681	=>	52350,
		6682	=>	52353,
		6683	=>	52355,
		6684	=>	52358,
		6685	=>	52360,
		6686	=>	52363,
		6687	=>	52365,
		6688	=>	52368,
		6689	=>	52370,
		6690	=>	52373,
		6691	=>	52375,
		6692	=>	52378,
		6693	=>	52380,
		6694	=>	52383,
		6695	=>	52385,
		6696	=>	52388,
		6697	=>	52390,
		6698	=>	52393,
		6699	=>	52395,
		6700	=>	52398,
		6701	=>	52400,
		6702	=>	52403,
		6703	=>	52405,
		6704	=>	52408,
		6705	=>	52411,
		6706	=>	52413,
		6707	=>	52416,
		6708	=>	52418,
		6709	=>	52421,
		6710	=>	52423,
		6711	=>	52426,
		6712	=>	52428,
		6713	=>	52431,
		6714	=>	52433,
		6715	=>	52436,
		6716	=>	52438,
		6717	=>	52441,
		6718	=>	52443,
		6719	=>	52446,
		6720	=>	52448,
		6721	=>	52451,
		6722	=>	52453,
		6723	=>	52456,
		6724	=>	52458,
		6725	=>	52461,
		6726	=>	52463,
		6727	=>	52466,
		6728	=>	52468,
		6729	=>	52471,
		6730	=>	52473,
		6731	=>	52476,
		6732	=>	52478,
		6733	=>	52481,
		6734	=>	52483,
		6735	=>	52486,
		6736	=>	52488,
		6737	=>	52491,
		6738	=>	52493,
		6739	=>	52496,
		6740	=>	52498,
		6741	=>	52501,
		6742	=>	52503,
		6743	=>	52506,
		6744	=>	52508,
		6745	=>	52511,
		6746	=>	52513,
		6747	=>	52516,
		6748	=>	52518,
		6749	=>	52521,
		6750	=>	52523,
		6751	=>	52526,
		6752	=>	52528,
		6753	=>	52531,
		6754	=>	52533,
		6755	=>	52536,
		6756	=>	52539,
		6757	=>	52541,
		6758	=>	52544,
		6759	=>	52546,
		6760	=>	52549,
		6761	=>	52551,
		6762	=>	52554,
		6763	=>	52556,
		6764	=>	52559,
		6765	=>	52561,
		6766	=>	52564,
		6767	=>	52566,
		6768	=>	52569,
		6769	=>	52571,
		6770	=>	52574,
		6771	=>	52576,
		6772	=>	52579,
		6773	=>	52581,
		6774	=>	52584,
		6775	=>	52586,
		6776	=>	52589,
		6777	=>	52591,
		6778	=>	52594,
		6779	=>	52596,
		6780	=>	52599,
		6781	=>	52601,
		6782	=>	52604,
		6783	=>	52606,
		6784	=>	52609,
		6785	=>	52611,
		6786	=>	52614,
		6787	=>	52616,
		6788	=>	52619,
		6789	=>	52621,
		6790	=>	52624,
		6791	=>	52626,
		6792	=>	52629,
		6793	=>	52631,
		6794	=>	52634,
		6795	=>	52636,
		6796	=>	52639,
		6797	=>	52641,
		6798	=>	52644,
		6799	=>	52646,
		6800	=>	52649,
		6801	=>	52651,
		6802	=>	52654,
		6803	=>	52656,
		6804	=>	52659,
		6805	=>	52661,
		6806	=>	52664,
		6807	=>	52666,
		6808	=>	52669,
		6809	=>	52671,
		6810	=>	52674,
		6811	=>	52676,
		6812	=>	52679,
		6813	=>	52681,
		6814	=>	52684,
		6815	=>	52686,
		6816	=>	52688,
		6817	=>	52691,
		6818	=>	52693,
		6819	=>	52696,
		6820	=>	52698,
		6821	=>	52701,
		6822	=>	52703,
		6823	=>	52706,
		6824	=>	52708,
		6825	=>	52711,
		6826	=>	52713,
		6827	=>	52716,
		6828	=>	52718,
		6829	=>	52721,
		6830	=>	52723,
		6831	=>	52726,
		6832	=>	52728,
		6833	=>	52731,
		6834	=>	52733,
		6835	=>	52736,
		6836	=>	52738,
		6837	=>	52741,
		6838	=>	52743,
		6839	=>	52746,
		6840	=>	52748,
		6841	=>	52751,
		6842	=>	52753,
		6843	=>	52756,
		6844	=>	52758,
		6845	=>	52761,
		6846	=>	52763,
		6847	=>	52766,
		6848	=>	52768,
		6849	=>	52771,
		6850	=>	52773,
		6851	=>	52776,
		6852	=>	52778,
		6853	=>	52781,
		6854	=>	52783,
		6855	=>	52786,
		6856	=>	52788,
		6857	=>	52791,
		6858	=>	52793,
		6859	=>	52796,
		6860	=>	52798,
		6861	=>	52801,
		6862	=>	52803,
		6863	=>	52806,
		6864	=>	52808,
		6865	=>	52810,
		6866	=>	52813,
		6867	=>	52815,
		6868	=>	52818,
		6869	=>	52820,
		6870	=>	52823,
		6871	=>	52825,
		6872	=>	52828,
		6873	=>	52830,
		6874	=>	52833,
		6875	=>	52835,
		6876	=>	52838,
		6877	=>	52840,
		6878	=>	52843,
		6879	=>	52845,
		6880	=>	52848,
		6881	=>	52850,
		6882	=>	52853,
		6883	=>	52855,
		6884	=>	52858,
		6885	=>	52860,
		6886	=>	52863,
		6887	=>	52865,
		6888	=>	52868,
		6889	=>	52870,
		6890	=>	52873,
		6891	=>	52875,
		6892	=>	52878,
		6893	=>	52880,
		6894	=>	52882,
		6895	=>	52885,
		6896	=>	52887,
		6897	=>	52890,
		6898	=>	52892,
		6899	=>	52895,
		6900	=>	52897,
		6901	=>	52900,
		6902	=>	52902,
		6903	=>	52905,
		6904	=>	52907,
		6905	=>	52910,
		6906	=>	52912,
		6907	=>	52915,
		6908	=>	52917,
		6909	=>	52920,
		6910	=>	52922,
		6911	=>	52925,
		6912	=>	52927,
		6913	=>	52930,
		6914	=>	52932,
		6915	=>	52935,
		6916	=>	52937,
		6917	=>	52939,
		6918	=>	52942,
		6919	=>	52944,
		6920	=>	52947,
		6921	=>	52949,
		6922	=>	52952,
		6923	=>	52954,
		6924	=>	52957,
		6925	=>	52959,
		6926	=>	52962,
		6927	=>	52964,
		6928	=>	52967,
		6929	=>	52969,
		6930	=>	52972,
		6931	=>	52974,
		6932	=>	52977,
		6933	=>	52979,
		6934	=>	52982,
		6935	=>	52984,
		6936	=>	52986,
		6937	=>	52989,
		6938	=>	52991,
		6939	=>	52994,
		6940	=>	52996,
		6941	=>	52999,
		6942	=>	53001,
		6943	=>	53004,
		6944	=>	53006,
		6945	=>	53009,
		6946	=>	53011,
		6947	=>	53014,
		6948	=>	53016,
		6949	=>	53019,
		6950	=>	53021,
		6951	=>	53024,
		6952	=>	53026,
		6953	=>	53028,
		6954	=>	53031,
		6955	=>	53033,
		6956	=>	53036,
		6957	=>	53038,
		6958	=>	53041,
		6959	=>	53043,
		6960	=>	53046,
		6961	=>	53048,
		6962	=>	53051,
		6963	=>	53053,
		6964	=>	53056,
		6965	=>	53058,
		6966	=>	53061,
		6967	=>	53063,
		6968	=>	53066,
		6969	=>	53068,
		6970	=>	53070,
		6971	=>	53073,
		6972	=>	53075,
		6973	=>	53078,
		6974	=>	53080,
		6975	=>	53083,
		6976	=>	53085,
		6977	=>	53088,
		6978	=>	53090,
		6979	=>	53093,
		6980	=>	53095,
		6981	=>	53098,
		6982	=>	53100,
		6983	=>	53102,
		6984	=>	53105,
		6985	=>	53107,
		6986	=>	53110,
		6987	=>	53112,
		6988	=>	53115,
		6989	=>	53117,
		6990	=>	53120,
		6991	=>	53122,
		6992	=>	53125,
		6993	=>	53127,
		6994	=>	53130,
		6995	=>	53132,
		6996	=>	53134,
		6997	=>	53137,
		6998	=>	53139,
		6999	=>	53142,
		7000	=>	53144,
		7001	=>	53147,
		7002	=>	53149,
		7003	=>	53152,
		7004	=>	53154,
		7005	=>	53157,
		7006	=>	53159,
		7007	=>	53162,
		7008	=>	53164,
		7009	=>	53166,
		7010	=>	53169,
		7011	=>	53171,
		7012	=>	53174,
		7013	=>	53176,
		7014	=>	53179,
		7015	=>	53181,
		7016	=>	53184,
		7017	=>	53186,
		7018	=>	53189,
		7019	=>	53191,
		7020	=>	53193,
		7021	=>	53196,
		7022	=>	53198,
		7023	=>	53201,
		7024	=>	53203,
		7025	=>	53206,
		7026	=>	53208,
		7027	=>	53211,
		7028	=>	53213,
		7029	=>	53216,
		7030	=>	53218,
		7031	=>	53221,
		7032	=>	53223,
		7033	=>	53225,
		7034	=>	53228,
		7035	=>	53230,
		7036	=>	53233,
		7037	=>	53235,
		7038	=>	53238,
		7039	=>	53240,
		7040	=>	53243,
		7041	=>	53245,
		7042	=>	53247,
		7043	=>	53250,
		7044	=>	53252,
		7045	=>	53255,
		7046	=>	53257,
		7047	=>	53260,
		7048	=>	53262,
		7049	=>	53265,
		7050	=>	53267,
		7051	=>	53270,
		7052	=>	53272,
		7053	=>	53274,
		7054	=>	53277,
		7055	=>	53279,
		7056	=>	53282,
		7057	=>	53284,
		7058	=>	53287,
		7059	=>	53289,
		7060	=>	53292,
		7061	=>	53294,
		7062	=>	53296,
		7063	=>	53299,
		7064	=>	53301,
		7065	=>	53304,
		7066	=>	53306,
		7067	=>	53309,
		7068	=>	53311,
		7069	=>	53314,
		7070	=>	53316,
		7071	=>	53319,
		7072	=>	53321,
		7073	=>	53323,
		7074	=>	53326,
		7075	=>	53328,
		7076	=>	53331,
		7077	=>	53333,
		7078	=>	53336,
		7079	=>	53338,
		7080	=>	53341,
		7081	=>	53343,
		7082	=>	53345,
		7083	=>	53348,
		7084	=>	53350,
		7085	=>	53353,
		7086	=>	53355,
		7087	=>	53358,
		7088	=>	53360,
		7089	=>	53363,
		7090	=>	53365,
		7091	=>	53367,
		7092	=>	53370,
		7093	=>	53372,
		7094	=>	53375,
		7095	=>	53377,
		7096	=>	53380,
		7097	=>	53382,
		7098	=>	53385,
		7099	=>	53387,
		7100	=>	53389,
		7101	=>	53392,
		7102	=>	53394,
		7103	=>	53397,
		7104	=>	53399,
		7105	=>	53402,
		7106	=>	53404,
		7107	=>	53406,
		7108	=>	53409,
		7109	=>	53411,
		7110	=>	53414,
		7111	=>	53416,
		7112	=>	53419,
		7113	=>	53421,
		7114	=>	53424,
		7115	=>	53426,
		7116	=>	53428,
		7117	=>	53431,
		7118	=>	53433,
		7119	=>	53436,
		7120	=>	53438,
		7121	=>	53441,
		7122	=>	53443,
		7123	=>	53446,
		7124	=>	53448,
		7125	=>	53450,
		7126	=>	53453,
		7127	=>	53455,
		7128	=>	53458,
		7129	=>	53460,
		7130	=>	53463,
		7131	=>	53465,
		7132	=>	53467,
		7133	=>	53470,
		7134	=>	53472,
		7135	=>	53475,
		7136	=>	53477,
		7137	=>	53480,
		7138	=>	53482,
		7139	=>	53484,
		7140	=>	53487,
		7141	=>	53489,
		7142	=>	53492,
		7143	=>	53494,
		7144	=>	53497,
		7145	=>	53499,
		7146	=>	53502,
		7147	=>	53504,
		7148	=>	53506,
		7149	=>	53509,
		7150	=>	53511,
		7151	=>	53514,
		7152	=>	53516,
		7153	=>	53519,
		7154	=>	53521,
		7155	=>	53523,
		7156	=>	53526,
		7157	=>	53528,
		7158	=>	53531,
		7159	=>	53533,
		7160	=>	53536,
		7161	=>	53538,
		7162	=>	53540,
		7163	=>	53543,
		7164	=>	53545,
		7165	=>	53548,
		7166	=>	53550,
		7167	=>	53553,
		7168	=>	53555,
		7169	=>	53557,
		7170	=>	53560,
		7171	=>	53562,
		7172	=>	53565,
		7173	=>	53567,
		7174	=>	53570,
		7175	=>	53572,
		7176	=>	53574,
		7177	=>	53577,
		7178	=>	53579,
		7179	=>	53582,
		7180	=>	53584,
		7181	=>	53587,
		7182	=>	53589,
		7183	=>	53591,
		7184	=>	53594,
		7185	=>	53596,
		7186	=>	53599,
		7187	=>	53601,
		7188	=>	53604,
		7189	=>	53606,
		7190	=>	53608,
		7191	=>	53611,
		7192	=>	53613,
		7193	=>	53616,
		7194	=>	53618,
		7195	=>	53620,
		7196	=>	53623,
		7197	=>	53625,
		7198	=>	53628,
		7199	=>	53630,
		7200	=>	53633,
		7201	=>	53635,
		7202	=>	53637,
		7203	=>	53640,
		7204	=>	53642,
		7205	=>	53645,
		7206	=>	53647,
		7207	=>	53650,
		7208	=>	53652,
		7209	=>	53654,
		7210	=>	53657,
		7211	=>	53659,
		7212	=>	53662,
		7213	=>	53664,
		7214	=>	53666,
		7215	=>	53669,
		7216	=>	53671,
		7217	=>	53674,
		7218	=>	53676,
		7219	=>	53679,
		7220	=>	53681,
		7221	=>	53683,
		7222	=>	53686,
		7223	=>	53688,
		7224	=>	53691,
		7225	=>	53693,
		7226	=>	53696,
		7227	=>	53698,
		7228	=>	53700,
		7229	=>	53703,
		7230	=>	53705,
		7231	=>	53708,
		7232	=>	53710,
		7233	=>	53712,
		7234	=>	53715,
		7235	=>	53717,
		7236	=>	53720,
		7237	=>	53722,
		7238	=>	53725,
		7239	=>	53727,
		7240	=>	53729,
		7241	=>	53732,
		7242	=>	53734,
		7243	=>	53737,
		7244	=>	53739,
		7245	=>	53741,
		7246	=>	53744,
		7247	=>	53746,
		7248	=>	53749,
		7249	=>	53751,
		7250	=>	53753,
		7251	=>	53756,
		7252	=>	53758,
		7253	=>	53761,
		7254	=>	53763,
		7255	=>	53766,
		7256	=>	53768,
		7257	=>	53770,
		7258	=>	53773,
		7259	=>	53775,
		7260	=>	53778,
		7261	=>	53780,
		7262	=>	53782,
		7263	=>	53785,
		7264	=>	53787,
		7265	=>	53790,
		7266	=>	53792,
		7267	=>	53794,
		7268	=>	53797,
		7269	=>	53799,
		7270	=>	53802,
		7271	=>	53804,
		7272	=>	53807,
		7273	=>	53809,
		7274	=>	53811,
		7275	=>	53814,
		7276	=>	53816,
		7277	=>	53819,
		7278	=>	53821,
		7279	=>	53823,
		7280	=>	53826,
		7281	=>	53828,
		7282	=>	53831,
		7283	=>	53833,
		7284	=>	53835,
		7285	=>	53838,
		7286	=>	53840,
		7287	=>	53843,
		7288	=>	53845,
		7289	=>	53847,
		7290	=>	53850,
		7291	=>	53852,
		7292	=>	53855,
		7293	=>	53857,
		7294	=>	53859,
		7295	=>	53862,
		7296	=>	53864,
		7297	=>	53867,
		7298	=>	53869,
		7299	=>	53871,
		7300	=>	53874,
		7301	=>	53876,
		7302	=>	53879,
		7303	=>	53881,
		7304	=>	53883,
		7305	=>	53886,
		7306	=>	53888,
		7307	=>	53891,
		7308	=>	53893,
		7309	=>	53895,
		7310	=>	53898,
		7311	=>	53900,
		7312	=>	53903,
		7313	=>	53905,
		7314	=>	53907,
		7315	=>	53910,
		7316	=>	53912,
		7317	=>	53915,
		7318	=>	53917,
		7319	=>	53919,
		7320	=>	53922,
		7321	=>	53924,
		7322	=>	53927,
		7323	=>	53929,
		7324	=>	53931,
		7325	=>	53934,
		7326	=>	53936,
		7327	=>	53939,
		7328	=>	53941,
		7329	=>	53943,
		7330	=>	53946,
		7331	=>	53948,
		7332	=>	53951,
		7333	=>	53953,
		7334	=>	53955,
		7335	=>	53958,
		7336	=>	53960,
		7337	=>	53963,
		7338	=>	53965,
		7339	=>	53967,
		7340	=>	53970,
		7341	=>	53972,
		7342	=>	53975,
		7343	=>	53977,
		7344	=>	53979,
		7345	=>	53982,
		7346	=>	53984,
		7347	=>	53987,
		7348	=>	53989,
		7349	=>	53991,
		7350	=>	53994,
		7351	=>	53996,
		7352	=>	53999,
		7353	=>	54001,
		7354	=>	54003,
		7355	=>	54006,
		7356	=>	54008,
		7357	=>	54011,
		7358	=>	54013,
		7359	=>	54015,
		7360	=>	54018,
		7361	=>	54020,
		7362	=>	54022,
		7363	=>	54025,
		7364	=>	54027,
		7365	=>	54030,
		7366	=>	54032,
		7367	=>	54034,
		7368	=>	54037,
		7369	=>	54039,
		7370	=>	54042,
		7371	=>	54044,
		7372	=>	54046,
		7373	=>	54049,
		7374	=>	54051,
		7375	=>	54054,
		7376	=>	54056,
		7377	=>	54058,
		7378	=>	54061,
		7379	=>	54063,
		7380	=>	54065,
		7381	=>	54068,
		7382	=>	54070,
		7383	=>	54073,
		7384	=>	54075,
		7385	=>	54077,
		7386	=>	54080,
		7387	=>	54082,
		7388	=>	54085,
		7389	=>	54087,
		7390	=>	54089,
		7391	=>	54092,
		7392	=>	54094,
		7393	=>	54097,
		7394	=>	54099,
		7395	=>	54101,
		7396	=>	54104,
		7397	=>	54106,
		7398	=>	54108,
		7399	=>	54111,
		7400	=>	54113,
		7401	=>	54116,
		7402	=>	54118,
		7403	=>	54120,
		7404	=>	54123,
		7405	=>	54125,
		7406	=>	54127,
		7407	=>	54130,
		7408	=>	54132,
		7409	=>	54135,
		7410	=>	54137,
		7411	=>	54139,
		7412	=>	54142,
		7413	=>	54144,
		7414	=>	54147,
		7415	=>	54149,
		7416	=>	54151,
		7417	=>	54154,
		7418	=>	54156,
		7419	=>	54158,
		7420	=>	54161,
		7421	=>	54163,
		7422	=>	54166,
		7423	=>	54168,
		7424	=>	54170,
		7425	=>	54173,
		7426	=>	54175,
		7427	=>	54177,
		7428	=>	54180,
		7429	=>	54182,
		7430	=>	54185,
		7431	=>	54187,
		7432	=>	54189,
		7433	=>	54192,
		7434	=>	54194,
		7435	=>	54196,
		7436	=>	54199,
		7437	=>	54201,
		7438	=>	54204,
		7439	=>	54206,
		7440	=>	54208,
		7441	=>	54211,
		7442	=>	54213,
		7443	=>	54216,
		7444	=>	54218,
		7445	=>	54220,
		7446	=>	54223,
		7447	=>	54225,
		7448	=>	54227,
		7449	=>	54230,
		7450	=>	54232,
		7451	=>	54234,
		7452	=>	54237,
		7453	=>	54239,
		7454	=>	54242,
		7455	=>	54244,
		7456	=>	54246,
		7457	=>	54249,
		7458	=>	54251,
		7459	=>	54253,
		7460	=>	54256,
		7461	=>	54258,
		7462	=>	54261,
		7463	=>	54263,
		7464	=>	54265,
		7465	=>	54268,
		7466	=>	54270,
		7467	=>	54272,
		7468	=>	54275,
		7469	=>	54277,
		7470	=>	54280,
		7471	=>	54282,
		7472	=>	54284,
		7473	=>	54287,
		7474	=>	54289,
		7475	=>	54291,
		7476	=>	54294,
		7477	=>	54296,
		7478	=>	54299,
		7479	=>	54301,
		7480	=>	54303,
		7481	=>	54306,
		7482	=>	54308,
		7483	=>	54310,
		7484	=>	54313,
		7485	=>	54315,
		7486	=>	54317,
		7487	=>	54320,
		7488	=>	54322,
		7489	=>	54325,
		7490	=>	54327,
		7491	=>	54329,
		7492	=>	54332,
		7493	=>	54334,
		7494	=>	54336,
		7495	=>	54339,
		7496	=>	54341,
		7497	=>	54343,
		7498	=>	54346,
		7499	=>	54348,
		7500	=>	54351,
		7501	=>	54353,
		7502	=>	54355,
		7503	=>	54358,
		7504	=>	54360,
		7505	=>	54362,
		7506	=>	54365,
		7507	=>	54367,
		7508	=>	54369,
		7509	=>	54372,
		7510	=>	54374,
		7511	=>	54377,
		7512	=>	54379,
		7513	=>	54381,
		7514	=>	54384,
		7515	=>	54386,
		7516	=>	54388,
		7517	=>	54391,
		7518	=>	54393,
		7519	=>	54395,
		7520	=>	54398,
		7521	=>	54400,
		7522	=>	54403,
		7523	=>	54405,
		7524	=>	54407,
		7525	=>	54410,
		7526	=>	54412,
		7527	=>	54414,
		7528	=>	54417,
		7529	=>	54419,
		7530	=>	54421,
		7531	=>	54424,
		7532	=>	54426,
		7533	=>	54428,
		7534	=>	54431,
		7535	=>	54433,
		7536	=>	54436,
		7537	=>	54438,
		7538	=>	54440,
		7539	=>	54443,
		7540	=>	54445,
		7541	=>	54447,
		7542	=>	54450,
		7543	=>	54452,
		7544	=>	54454,
		7545	=>	54457,
		7546	=>	54459,
		7547	=>	54461,
		7548	=>	54464,
		7549	=>	54466,
		7550	=>	54469,
		7551	=>	54471,
		7552	=>	54473,
		7553	=>	54476,
		7554	=>	54478,
		7555	=>	54480,
		7556	=>	54483,
		7557	=>	54485,
		7558	=>	54487,
		7559	=>	54490,
		7560	=>	54492,
		7561	=>	54494,
		7562	=>	54497,
		7563	=>	54499,
		7564	=>	54501,
		7565	=>	54504,
		7566	=>	54506,
		7567	=>	54508,
		7568	=>	54511,
		7569	=>	54513,
		7570	=>	54516,
		7571	=>	54518,
		7572	=>	54520,
		7573	=>	54523,
		7574	=>	54525,
		7575	=>	54527,
		7576	=>	54530,
		7577	=>	54532,
		7578	=>	54534,
		7579	=>	54537,
		7580	=>	54539,
		7581	=>	54541,
		7582	=>	54544,
		7583	=>	54546,
		7584	=>	54548,
		7585	=>	54551,
		7586	=>	54553,
		7587	=>	54555,
		7588	=>	54558,
		7589	=>	54560,
		7590	=>	54562,
		7591	=>	54565,
		7592	=>	54567,
		7593	=>	54570,
		7594	=>	54572,
		7595	=>	54574,
		7596	=>	54577,
		7597	=>	54579,
		7598	=>	54581,
		7599	=>	54584,
		7600	=>	54586,
		7601	=>	54588,
		7602	=>	54591,
		7603	=>	54593,
		7604	=>	54595,
		7605	=>	54598,
		7606	=>	54600,
		7607	=>	54602,
		7608	=>	54605,
		7609	=>	54607,
		7610	=>	54609,
		7611	=>	54612,
		7612	=>	54614,
		7613	=>	54616,
		7614	=>	54619,
		7615	=>	54621,
		7616	=>	54623,
		7617	=>	54626,
		7618	=>	54628,
		7619	=>	54630,
		7620	=>	54633,
		7621	=>	54635,
		7622	=>	54637,
		7623	=>	54640,
		7624	=>	54642,
		7625	=>	54644,
		7626	=>	54647,
		7627	=>	54649,
		7628	=>	54651,
		7629	=>	54654,
		7630	=>	54656,
		7631	=>	54659,
		7632	=>	54661,
		7633	=>	54663,
		7634	=>	54666,
		7635	=>	54668,
		7636	=>	54670,
		7637	=>	54673,
		7638	=>	54675,
		7639	=>	54677,
		7640	=>	54680,
		7641	=>	54682,
		7642	=>	54684,
		7643	=>	54687,
		7644	=>	54689,
		7645	=>	54691,
		7646	=>	54694,
		7647	=>	54696,
		7648	=>	54698,
		7649	=>	54701,
		7650	=>	54703,
		7651	=>	54705,
		7652	=>	54708,
		7653	=>	54710,
		7654	=>	54712,
		7655	=>	54715,
		7656	=>	54717,
		7657	=>	54719,
		7658	=>	54722,
		7659	=>	54724,
		7660	=>	54726,
		7661	=>	54729,
		7662	=>	54731,
		7663	=>	54733,
		7664	=>	54736,
		7665	=>	54738,
		7666	=>	54740,
		7667	=>	54743,
		7668	=>	54745,
		7669	=>	54747,
		7670	=>	54750,
		7671	=>	54752,
		7672	=>	54754,
		7673	=>	54757,
		7674	=>	54759,
		7675	=>	54761,
		7676	=>	54763,
		7677	=>	54766,
		7678	=>	54768,
		7679	=>	54770,
		7680	=>	54773,
		7681	=>	54775,
		7682	=>	54777,
		7683	=>	54780,
		7684	=>	54782,
		7685	=>	54784,
		7686	=>	54787,
		7687	=>	54789,
		7688	=>	54791,
		7689	=>	54794,
		7690	=>	54796,
		7691	=>	54798,
		7692	=>	54801,
		7693	=>	54803,
		7694	=>	54805,
		7695	=>	54808,
		7696	=>	54810,
		7697	=>	54812,
		7698	=>	54815,
		7699	=>	54817,
		7700	=>	54819,
		7701	=>	54822,
		7702	=>	54824,
		7703	=>	54826,
		7704	=>	54829,
		7705	=>	54831,
		7706	=>	54833,
		7707	=>	54836,
		7708	=>	54838,
		7709	=>	54840,
		7710	=>	54843,
		7711	=>	54845,
		7712	=>	54847,
		7713	=>	54850,
		7714	=>	54852,
		7715	=>	54854,
		7716	=>	54856,
		7717	=>	54859,
		7718	=>	54861,
		7719	=>	54863,
		7720	=>	54866,
		7721	=>	54868,
		7722	=>	54870,
		7723	=>	54873,
		7724	=>	54875,
		7725	=>	54877,
		7726	=>	54880,
		7727	=>	54882,
		7728	=>	54884,
		7729	=>	54887,
		7730	=>	54889,
		7731	=>	54891,
		7732	=>	54894,
		7733	=>	54896,
		7734	=>	54898,
		7735	=>	54901,
		7736	=>	54903,
		7737	=>	54905,
		7738	=>	54907,
		7739	=>	54910,
		7740	=>	54912,
		7741	=>	54914,
		7742	=>	54917,
		7743	=>	54919,
		7744	=>	54921,
		7745	=>	54924,
		7746	=>	54926,
		7747	=>	54928,
		7748	=>	54931,
		7749	=>	54933,
		7750	=>	54935,
		7751	=>	54938,
		7752	=>	54940,
		7753	=>	54942,
		7754	=>	54945,
		7755	=>	54947,
		7756	=>	54949,
		7757	=>	54951,
		7758	=>	54954,
		7759	=>	54956,
		7760	=>	54958,
		7761	=>	54961,
		7762	=>	54963,
		7763	=>	54965,
		7764	=>	54968,
		7765	=>	54970,
		7766	=>	54972,
		7767	=>	54975,
		7768	=>	54977,
		7769	=>	54979,
		7770	=>	54981,
		7771	=>	54984,
		7772	=>	54986,
		7773	=>	54988,
		7774	=>	54991,
		7775	=>	54993,
		7776	=>	54995,
		7777	=>	54998,
		7778	=>	55000,
		7779	=>	55002,
		7780	=>	55005,
		7781	=>	55007,
		7782	=>	55009,
		7783	=>	55011,
		7784	=>	55014,
		7785	=>	55016,
		7786	=>	55018,
		7787	=>	55021,
		7788	=>	55023,
		7789	=>	55025,
		7790	=>	55028,
		7791	=>	55030,
		7792	=>	55032,
		7793	=>	55035,
		7794	=>	55037,
		7795	=>	55039,
		7796	=>	55041,
		7797	=>	55044,
		7798	=>	55046,
		7799	=>	55048,
		7800	=>	55051,
		7801	=>	55053,
		7802	=>	55055,
		7803	=>	55058,
		7804	=>	55060,
		7805	=>	55062,
		7806	=>	55064,
		7807	=>	55067,
		7808	=>	55069,
		7809	=>	55071,
		7810	=>	55074,
		7811	=>	55076,
		7812	=>	55078,
		7813	=>	55081,
		7814	=>	55083,
		7815	=>	55085,
		7816	=>	55087,
		7817	=>	55090,
		7818	=>	55092,
		7819	=>	55094,
		7820	=>	55097,
		7821	=>	55099,
		7822	=>	55101,
		7823	=>	55104,
		7824	=>	55106,
		7825	=>	55108,
		7826	=>	55110,
		7827	=>	55113,
		7828	=>	55115,
		7829	=>	55117,
		7830	=>	55120,
		7831	=>	55122,
		7832	=>	55124,
		7833	=>	55127,
		7834	=>	55129,
		7835	=>	55131,
		7836	=>	55133,
		7837	=>	55136,
		7838	=>	55138,
		7839	=>	55140,
		7840	=>	55143,
		7841	=>	55145,
		7842	=>	55147,
		7843	=>	55150,
		7844	=>	55152,
		7845	=>	55154,
		7846	=>	55156,
		7847	=>	55159,
		7848	=>	55161,
		7849	=>	55163,
		7850	=>	55166,
		7851	=>	55168,
		7852	=>	55170,
		7853	=>	55172,
		7854	=>	55175,
		7855	=>	55177,
		7856	=>	55179,
		7857	=>	55182,
		7858	=>	55184,
		7859	=>	55186,
		7860	=>	55189,
		7861	=>	55191,
		7862	=>	55193,
		7863	=>	55195,
		7864	=>	55198,
		7865	=>	55200,
		7866	=>	55202,
		7867	=>	55205,
		7868	=>	55207,
		7869	=>	55209,
		7870	=>	55211,
		7871	=>	55214,
		7872	=>	55216,
		7873	=>	55218,
		7874	=>	55221,
		7875	=>	55223,
		7876	=>	55225,
		7877	=>	55227,
		7878	=>	55230,
		7879	=>	55232,
		7880	=>	55234,
		7881	=>	55237,
		7882	=>	55239,
		7883	=>	55241,
		7884	=>	55243,
		7885	=>	55246,
		7886	=>	55248,
		7887	=>	55250,
		7888	=>	55253,
		7889	=>	55255,
		7890	=>	55257,
		7891	=>	55259,
		7892	=>	55262,
		7893	=>	55264,
		7894	=>	55266,
		7895	=>	55269,
		7896	=>	55271,
		7897	=>	55273,
		7898	=>	55275,
		7899	=>	55278,
		7900	=>	55280,
		7901	=>	55282,
		7902	=>	55285,
		7903	=>	55287,
		7904	=>	55289,
		7905	=>	55291,
		7906	=>	55294,
		7907	=>	55296,
		7908	=>	55298,
		7909	=>	55301,
		7910	=>	55303,
		7911	=>	55305,
		7912	=>	55307,
		7913	=>	55310,
		7914	=>	55312,
		7915	=>	55314,
		7916	=>	55316,
		7917	=>	55319,
		7918	=>	55321,
		7919	=>	55323,
		7920	=>	55326,
		7921	=>	55328,
		7922	=>	55330,
		7923	=>	55332,
		7924	=>	55335,
		7925	=>	55337,
		7926	=>	55339,
		7927	=>	55342,
		7928	=>	55344,
		7929	=>	55346,
		7930	=>	55348,
		7931	=>	55351,
		7932	=>	55353,
		7933	=>	55355,
		7934	=>	55357,
		7935	=>	55360,
		7936	=>	55362,
		7937	=>	55364,
		7938	=>	55367,
		7939	=>	55369,
		7940	=>	55371,
		7941	=>	55373,
		7942	=>	55376,
		7943	=>	55378,
		7944	=>	55380,
		7945	=>	55382,
		7946	=>	55385,
		7947	=>	55387,
		7948	=>	55389,
		7949	=>	55392,
		7950	=>	55394,
		7951	=>	55396,
		7952	=>	55398,
		7953	=>	55401,
		7954	=>	55403,
		7955	=>	55405,
		7956	=>	55407,
		7957	=>	55410,
		7958	=>	55412,
		7959	=>	55414,
		7960	=>	55417,
		7961	=>	55419,
		7962	=>	55421,
		7963	=>	55423,
		7964	=>	55426,
		7965	=>	55428,
		7966	=>	55430,
		7967	=>	55432,
		7968	=>	55435,
		7969	=>	55437,
		7970	=>	55439,
		7971	=>	55442,
		7972	=>	55444,
		7973	=>	55446,
		7974	=>	55448,
		7975	=>	55451,
		7976	=>	55453,
		7977	=>	55455,
		7978	=>	55457,
		7979	=>	55460,
		7980	=>	55462,
		7981	=>	55464,
		7982	=>	55466,
		7983	=>	55469,
		7984	=>	55471,
		7985	=>	55473,
		7986	=>	55476,
		7987	=>	55478,
		7988	=>	55480,
		7989	=>	55482,
		7990	=>	55485,
		7991	=>	55487,
		7992	=>	55489,
		7993	=>	55491,
		7994	=>	55494,
		7995	=>	55496,
		7996	=>	55498,
		7997	=>	55500,
		7998	=>	55503,
		7999	=>	55505,
		8000	=>	55507,
		8001	=>	55509,
		8002	=>	55512,
		8003	=>	55514,
		8004	=>	55516,
		8005	=>	55519,
		8006	=>	55521,
		8007	=>	55523,
		8008	=>	55525,
		8009	=>	55528,
		8010	=>	55530,
		8011	=>	55532,
		8012	=>	55534,
		8013	=>	55537,
		8014	=>	55539,
		8015	=>	55541,
		8016	=>	55543,
		8017	=>	55546,
		8018	=>	55548,
		8019	=>	55550,
		8020	=>	55552,
		8021	=>	55555,
		8022	=>	55557,
		8023	=>	55559,
		8024	=>	55561,
		8025	=>	55564,
		8026	=>	55566,
		8027	=>	55568,
		8028	=>	55570,
		8029	=>	55573,
		8030	=>	55575,
		8031	=>	55577,
		8032	=>	55579,
		8033	=>	55582,
		8034	=>	55584,
		8035	=>	55586,
		8036	=>	55589,
		8037	=>	55591,
		8038	=>	55593,
		8039	=>	55595,
		8040	=>	55598,
		8041	=>	55600,
		8042	=>	55602,
		8043	=>	55604,
		8044	=>	55607,
		8045	=>	55609,
		8046	=>	55611,
		8047	=>	55613,
		8048	=>	55616,
		8049	=>	55618,
		8050	=>	55620,
		8051	=>	55622,
		8052	=>	55625,
		8053	=>	55627,
		8054	=>	55629,
		8055	=>	55631,
		8056	=>	55634,
		8057	=>	55636,
		8058	=>	55638,
		8059	=>	55640,
		8060	=>	55643,
		8061	=>	55645,
		8062	=>	55647,
		8063	=>	55649,
		8064	=>	55652,
		8065	=>	55654,
		8066	=>	55656,
		8067	=>	55658,
		8068	=>	55661,
		8069	=>	55663,
		8070	=>	55665,
		8071	=>	55667,
		8072	=>	55670,
		8073	=>	55672,
		8074	=>	55674,
		8075	=>	55676,
		8076	=>	55679,
		8077	=>	55681,
		8078	=>	55683,
		8079	=>	55685,
		8080	=>	55687,
		8081	=>	55690,
		8082	=>	55692,
		8083	=>	55694,
		8084	=>	55696,
		8085	=>	55699,
		8086	=>	55701,
		8087	=>	55703,
		8088	=>	55705,
		8089	=>	55708,
		8090	=>	55710,
		8091	=>	55712,
		8092	=>	55714,
		8093	=>	55717,
		8094	=>	55719,
		8095	=>	55721,
		8096	=>	55723,
		8097	=>	55726,
		8098	=>	55728,
		8099	=>	55730,
		8100	=>	55732,
		8101	=>	55735,
		8102	=>	55737,
		8103	=>	55739,
		8104	=>	55741,
		8105	=>	55744,
		8106	=>	55746,
		8107	=>	55748,
		8108	=>	55750,
		8109	=>	55753,
		8110	=>	55755,
		8111	=>	55757,
		8112	=>	55759,
		8113	=>	55761,
		8114	=>	55764,
		8115	=>	55766,
		8116	=>	55768,
		8117	=>	55770,
		8118	=>	55773,
		8119	=>	55775,
		8120	=>	55777,
		8121	=>	55779,
		8122	=>	55782,
		8123	=>	55784,
		8124	=>	55786,
		8125	=>	55788,
		8126	=>	55791,
		8127	=>	55793,
		8128	=>	55795,
		8129	=>	55797,
		8130	=>	55799,
		8131	=>	55802,
		8132	=>	55804,
		8133	=>	55806,
		8134	=>	55808,
		8135	=>	55811,
		8136	=>	55813,
		8137	=>	55815,
		8138	=>	55817,
		8139	=>	55820,
		8140	=>	55822,
		8141	=>	55824,
		8142	=>	55826,
		8143	=>	55829,
		8144	=>	55831,
		8145	=>	55833,
		8146	=>	55835,
		8147	=>	55837,
		8148	=>	55840,
		8149	=>	55842,
		8150	=>	55844,
		8151	=>	55846,
		8152	=>	55849,
		8153	=>	55851,
		8154	=>	55853,
		8155	=>	55855,
		8156	=>	55858,
		8157	=>	55860,
		8158	=>	55862,
		8159	=>	55864,
		8160	=>	55866,
		8161	=>	55869,
		8162	=>	55871,
		8163	=>	55873,
		8164	=>	55875,
		8165	=>	55878,
		8166	=>	55880,
		8167	=>	55882,
		8168	=>	55884,
		8169	=>	55886,
		8170	=>	55889,
		8171	=>	55891,
		8172	=>	55893,
		8173	=>	55895,
		8174	=>	55898,
		8175	=>	55900,
		8176	=>	55902,
		8177	=>	55904,
		8178	=>	55907,
		8179	=>	55909,
		8180	=>	55911,
		8181	=>	55913,
		8182	=>	55915,
		8183	=>	55918,
		8184	=>	55920,
		8185	=>	55922,
		8186	=>	55924,
		8187	=>	55927,
		8188	=>	55929,
		8189	=>	55931,
		8190	=>	55933,
		8191	=>	55935,
		8192	=>	55938,
		8193	=>	55940,
		8194	=>	55942,
		8195	=>	55944,
		8196	=>	55947,
		8197	=>	55949,
		8198	=>	55951,
		8199	=>	55953,
		8200	=>	55955,
		8201	=>	55958,
		8202	=>	55960,
		8203	=>	55962,
		8204	=>	55964,
		8205	=>	55966,
		8206	=>	55969,
		8207	=>	55971,
		8208	=>	55973,
		8209	=>	55975,
		8210	=>	55978,
		8211	=>	55980,
		8212	=>	55982,
		8213	=>	55984,
		8214	=>	55986,
		8215	=>	55989,
		8216	=>	55991,
		8217	=>	55993,
		8218	=>	55995,
		8219	=>	55998,
		8220	=>	56000,
		8221	=>	56002,
		8222	=>	56004,
		8223	=>	56006,
		8224	=>	56009,
		8225	=>	56011,
		8226	=>	56013,
		8227	=>	56015,
		8228	=>	56017,
		8229	=>	56020,
		8230	=>	56022,
		8231	=>	56024,
		8232	=>	56026,
		8233	=>	56029,
		8234	=>	56031,
		8235	=>	56033,
		8236	=>	56035,
		8237	=>	56037,
		8238	=>	56040,
		8239	=>	56042,
		8240	=>	56044,
		8241	=>	56046,
		8242	=>	56048,
		8243	=>	56051,
		8244	=>	56053,
		8245	=>	56055,
		8246	=>	56057,
		8247	=>	56059,
		8248	=>	56062,
		8249	=>	56064,
		8250	=>	56066,
		8251	=>	56068,
		8252	=>	56071,
		8253	=>	56073,
		8254	=>	56075,
		8255	=>	56077,
		8256	=>	56079,
		8257	=>	56082,
		8258	=>	56084,
		8259	=>	56086,
		8260	=>	56088,
		8261	=>	56090,
		8262	=>	56093,
		8263	=>	56095,
		8264	=>	56097,
		8265	=>	56099,
		8266	=>	56101,
		8267	=>	56104,
		8268	=>	56106,
		8269	=>	56108,
		8270	=>	56110,
		8271	=>	56112,
		8272	=>	56115,
		8273	=>	56117,
		8274	=>	56119,
		8275	=>	56121,
		8276	=>	56123,
		8277	=>	56126,
		8278	=>	56128,
		8279	=>	56130,
		8280	=>	56132,
		8281	=>	56134,
		8282	=>	56137,
		8283	=>	56139,
		8284	=>	56141,
		8285	=>	56143,
		8286	=>	56145,
		8287	=>	56148,
		8288	=>	56150,
		8289	=>	56152,
		8290	=>	56154,
		8291	=>	56156,
		8292	=>	56159,
		8293	=>	56161,
		8294	=>	56163,
		8295	=>	56165,
		8296	=>	56167,
		8297	=>	56170,
		8298	=>	56172,
		8299	=>	56174,
		8300	=>	56176,
		8301	=>	56178,
		8302	=>	56181,
		8303	=>	56183,
		8304	=>	56185,
		8305	=>	56187,
		8306	=>	56189,
		8307	=>	56192,
		8308	=>	56194,
		8309	=>	56196,
		8310	=>	56198,
		8311	=>	56200,
		8312	=>	56203,
		8313	=>	56205,
		8314	=>	56207,
		8315	=>	56209,
		8316	=>	56211,
		8317	=>	56214,
		8318	=>	56216,
		8319	=>	56218,
		8320	=>	56220,
		8321	=>	56222,
		8322	=>	56225,
		8323	=>	56227,
		8324	=>	56229,
		8325	=>	56231,
		8326	=>	56233,
		8327	=>	56236,
		8328	=>	56238,
		8329	=>	56240,
		8330	=>	56242,
		8331	=>	56244,
		8332	=>	56247,
		8333	=>	56249,
		8334	=>	56251,
		8335	=>	56253,
		8336	=>	56255,
		8337	=>	56257,
		8338	=>	56260,
		8339	=>	56262,
		8340	=>	56264,
		8341	=>	56266,
		8342	=>	56268,
		8343	=>	56271,
		8344	=>	56273,
		8345	=>	56275,
		8346	=>	56277,
		8347	=>	56279,
		8348	=>	56282,
		8349	=>	56284,
		8350	=>	56286,
		8351	=>	56288,
		8352	=>	56290,
		8353	=>	56292,
		8354	=>	56295,
		8355	=>	56297,
		8356	=>	56299,
		8357	=>	56301,
		8358	=>	56303,
		8359	=>	56306,
		8360	=>	56308,
		8361	=>	56310,
		8362	=>	56312,
		8363	=>	56314,
		8364	=>	56317,
		8365	=>	56319,
		8366	=>	56321,
		8367	=>	56323,
		8368	=>	56325,
		8369	=>	56327,
		8370	=>	56330,
		8371	=>	56332,
		8372	=>	56334,
		8373	=>	56336,
		8374	=>	56338,
		8375	=>	56341,
		8376	=>	56343,
		8377	=>	56345,
		8378	=>	56347,
		8379	=>	56349,
		8380	=>	56351,
		8381	=>	56354,
		8382	=>	56356,
		8383	=>	56358,
		8384	=>	56360,
		8385	=>	56362,
		8386	=>	56365,
		8387	=>	56367,
		8388	=>	56369,
		8389	=>	56371,
		8390	=>	56373,
		8391	=>	56375,
		8392	=>	56378,
		8393	=>	56380,
		8394	=>	56382,
		8395	=>	56384,
		8396	=>	56386,
		8397	=>	56389,
		8398	=>	56391,
		8399	=>	56393,
		8400	=>	56395,
		8401	=>	56397,
		8402	=>	56399,
		8403	=>	56402,
		8404	=>	56404,
		8405	=>	56406,
		8406	=>	56408,
		8407	=>	56410,
		8408	=>	56412,
		8409	=>	56415,
		8410	=>	56417,
		8411	=>	56419,
		8412	=>	56421,
		8413	=>	56423,
		8414	=>	56425,
		8415	=>	56428,
		8416	=>	56430,
		8417	=>	56432,
		8418	=>	56434,
		8419	=>	56436,
		8420	=>	56439,
		8421	=>	56441,
		8422	=>	56443,
		8423	=>	56445,
		8424	=>	56447,
		8425	=>	56449,
		8426	=>	56452,
		8427	=>	56454,
		8428	=>	56456,
		8429	=>	56458,
		8430	=>	56460,
		8431	=>	56462,
		8432	=>	56465,
		8433	=>	56467,
		8434	=>	56469,
		8435	=>	56471,
		8436	=>	56473,
		8437	=>	56475,
		8438	=>	56478,
		8439	=>	56480,
		8440	=>	56482,
		8441	=>	56484,
		8442	=>	56486,
		8443	=>	56488,
		8444	=>	56491,
		8445	=>	56493,
		8446	=>	56495,
		8447	=>	56497,
		8448	=>	56499,
		8449	=>	56501,
		8450	=>	56504,
		8451	=>	56506,
		8452	=>	56508,
		8453	=>	56510,
		8454	=>	56512,
		8455	=>	56514,
		8456	=>	56517,
		8457	=>	56519,
		8458	=>	56521,
		8459	=>	56523,
		8460	=>	56525,
		8461	=>	56527,
		8462	=>	56530,
		8463	=>	56532,
		8464	=>	56534,
		8465	=>	56536,
		8466	=>	56538,
		8467	=>	56540,
		8468	=>	56543,
		8469	=>	56545,
		8470	=>	56547,
		8471	=>	56549,
		8472	=>	56551,
		8473	=>	56553,
		8474	=>	56556,
		8475	=>	56558,
		8476	=>	56560,
		8477	=>	56562,
		8478	=>	56564,
		8479	=>	56566,
		8480	=>	56568,
		8481	=>	56571,
		8482	=>	56573,
		8483	=>	56575,
		8484	=>	56577,
		8485	=>	56579,
		8486	=>	56581,
		8487	=>	56584,
		8488	=>	56586,
		8489	=>	56588,
		8490	=>	56590,
		8491	=>	56592,
		8492	=>	56594,
		8493	=>	56597,
		8494	=>	56599,
		8495	=>	56601,
		8496	=>	56603,
		8497	=>	56605,
		8498	=>	56607,
		8499	=>	56609,
		8500	=>	56612,
		8501	=>	56614,
		8502	=>	56616,
		8503	=>	56618,
		8504	=>	56620,
		8505	=>	56622,
		8506	=>	56625,
		8507	=>	56627,
		8508	=>	56629,
		8509	=>	56631,
		8510	=>	56633,
		8511	=>	56635,
		8512	=>	56637,
		8513	=>	56640,
		8514	=>	56642,
		8515	=>	56644,
		8516	=>	56646,
		8517	=>	56648,
		8518	=>	56650,
		8519	=>	56653,
		8520	=>	56655,
		8521	=>	56657,
		8522	=>	56659,
		8523	=>	56661,
		8524	=>	56663,
		8525	=>	56665,
		8526	=>	56668,
		8527	=>	56670,
		8528	=>	56672,
		8529	=>	56674,
		8530	=>	56676,
		8531	=>	56678,
		8532	=>	56680,
		8533	=>	56683,
		8534	=>	56685,
		8535	=>	56687,
		8536	=>	56689,
		8537	=>	56691,
		8538	=>	56693,
		8539	=>	56695,
		8540	=>	56698,
		8541	=>	56700,
		8542	=>	56702,
		8543	=>	56704,
		8544	=>	56706,
		8545	=>	56708,
		8546	=>	56711,
		8547	=>	56713,
		8548	=>	56715,
		8549	=>	56717,
		8550	=>	56719,
		8551	=>	56721,
		8552	=>	56723,
		8553	=>	56726,
		8554	=>	56728,
		8555	=>	56730,
		8556	=>	56732,
		8557	=>	56734,
		8558	=>	56736,
		8559	=>	56738,
		8560	=>	56741,
		8561	=>	56743,
		8562	=>	56745,
		8563	=>	56747,
		8564	=>	56749,
		8565	=>	56751,
		8566	=>	56753,
		8567	=>	56755,
		8568	=>	56758,
		8569	=>	56760,
		8570	=>	56762,
		8571	=>	56764,
		8572	=>	56766,
		8573	=>	56768,
		8574	=>	56770,
		8575	=>	56773,
		8576	=>	56775,
		8577	=>	56777,
		8578	=>	56779,
		8579	=>	56781,
		8580	=>	56783,
		8581	=>	56785,
		8582	=>	56788,
		8583	=>	56790,
		8584	=>	56792,
		8585	=>	56794,
		8586	=>	56796,
		8587	=>	56798,
		8588	=>	56800,
		8589	=>	56803,
		8590	=>	56805,
		8591	=>	56807,
		8592	=>	56809,
		8593	=>	56811,
		8594	=>	56813,
		8595	=>	56815,
		8596	=>	56817,
		8597	=>	56820,
		8598	=>	56822,
		8599	=>	56824,
		8600	=>	56826,
		8601	=>	56828,
		8602	=>	56830,
		8603	=>	56832,
		8604	=>	56835,
		8605	=>	56837,
		8606	=>	56839,
		8607	=>	56841,
		8608	=>	56843,
		8609	=>	56845,
		8610	=>	56847,
		8611	=>	56849,
		8612	=>	56852,
		8613	=>	56854,
		8614	=>	56856,
		8615	=>	56858,
		8616	=>	56860,
		8617	=>	56862,
		8618	=>	56864,
		8619	=>	56866,
		8620	=>	56869,
		8621	=>	56871,
		8622	=>	56873,
		8623	=>	56875,
		8624	=>	56877,
		8625	=>	56879,
		8626	=>	56881,
		8627	=>	56884,
		8628	=>	56886,
		8629	=>	56888,
		8630	=>	56890,
		8631	=>	56892,
		8632	=>	56894,
		8633	=>	56896,
		8634	=>	56898,
		8635	=>	56901,
		8636	=>	56903,
		8637	=>	56905,
		8638	=>	56907,
		8639	=>	56909,
		8640	=>	56911,
		8641	=>	56913,
		8642	=>	56915,
		8643	=>	56918,
		8644	=>	56920,
		8645	=>	56922,
		8646	=>	56924,
		8647	=>	56926,
		8648	=>	56928,
		8649	=>	56930,
		8650	=>	56932,
		8651	=>	56934,
		8652	=>	56937,
		8653	=>	56939,
		8654	=>	56941,
		8655	=>	56943,
		8656	=>	56945,
		8657	=>	56947,
		8658	=>	56949,
		8659	=>	56951,
		8660	=>	56954,
		8661	=>	56956,
		8662	=>	56958,
		8663	=>	56960,
		8664	=>	56962,
		8665	=>	56964,
		8666	=>	56966,
		8667	=>	56968,
		8668	=>	56971,
		8669	=>	56973,
		8670	=>	56975,
		8671	=>	56977,
		8672	=>	56979,
		8673	=>	56981,
		8674	=>	56983,
		8675	=>	56985,
		8676	=>	56987,
		8677	=>	56990,
		8678	=>	56992,
		8679	=>	56994,
		8680	=>	56996,
		8681	=>	56998,
		8682	=>	57000,
		8683	=>	57002,
		8684	=>	57004,
		8685	=>	57006,
		8686	=>	57009,
		8687	=>	57011,
		8688	=>	57013,
		8689	=>	57015,
		8690	=>	57017,
		8691	=>	57019,
		8692	=>	57021,
		8693	=>	57023,
		8694	=>	57026,
		8695	=>	57028,
		8696	=>	57030,
		8697	=>	57032,
		8698	=>	57034,
		8699	=>	57036,
		8700	=>	57038,
		8701	=>	57040,
		8702	=>	57042,
		8703	=>	57045,
		8704	=>	57047,
		8705	=>	57049,
		8706	=>	57051,
		8707	=>	57053,
		8708	=>	57055,
		8709	=>	57057,
		8710	=>	57059,
		8711	=>	57061,
		8712	=>	57063,
		8713	=>	57066,
		8714	=>	57068,
		8715	=>	57070,
		8716	=>	57072,
		8717	=>	57074,
		8718	=>	57076,
		8719	=>	57078,
		8720	=>	57080,
		8721	=>	57082,
		8722	=>	57085,
		8723	=>	57087,
		8724	=>	57089,
		8725	=>	57091,
		8726	=>	57093,
		8727	=>	57095,
		8728	=>	57097,
		8729	=>	57099,
		8730	=>	57101,
		8731	=>	57103,
		8732	=>	57106,
		8733	=>	57108,
		8734	=>	57110,
		8735	=>	57112,
		8736	=>	57114,
		8737	=>	57116,
		8738	=>	57118,
		8739	=>	57120,
		8740	=>	57122,
		8741	=>	57125,
		8742	=>	57127,
		8743	=>	57129,
		8744	=>	57131,
		8745	=>	57133,
		8746	=>	57135,
		8747	=>	57137,
		8748	=>	57139,
		8749	=>	57141,
		8750	=>	57143,
		8751	=>	57146,
		8752	=>	57148,
		8753	=>	57150,
		8754	=>	57152,
		8755	=>	57154,
		8756	=>	57156,
		8757	=>	57158,
		8758	=>	57160,
		8759	=>	57162,
		8760	=>	57164,
		8761	=>	57167,
		8762	=>	57169,
		8763	=>	57171,
		8764	=>	57173,
		8765	=>	57175,
		8766	=>	57177,
		8767	=>	57179,
		8768	=>	57181,
		8769	=>	57183,
		8770	=>	57185,
		8771	=>	57187,
		8772	=>	57190,
		8773	=>	57192,
		8774	=>	57194,
		8775	=>	57196,
		8776	=>	57198,
		8777	=>	57200,
		8778	=>	57202,
		8779	=>	57204,
		8780	=>	57206,
		8781	=>	57208,
		8782	=>	57210,
		8783	=>	57213,
		8784	=>	57215,
		8785	=>	57217,
		8786	=>	57219,
		8787	=>	57221,
		8788	=>	57223,
		8789	=>	57225,
		8790	=>	57227,
		8791	=>	57229,
		8792	=>	57231,
		8793	=>	57233,
		8794	=>	57236,
		8795	=>	57238,
		8796	=>	57240,
		8797	=>	57242,
		8798	=>	57244,
		8799	=>	57246,
		8800	=>	57248,
		8801	=>	57250,
		8802	=>	57252,
		8803	=>	57254,
		8804	=>	57256,
		8805	=>	57259,
		8806	=>	57261,
		8807	=>	57263,
		8808	=>	57265,
		8809	=>	57267,
		8810	=>	57269,
		8811	=>	57271,
		8812	=>	57273,
		8813	=>	57275,
		8814	=>	57277,
		8815	=>	57279,
		8816	=>	57282,
		8817	=>	57284,
		8818	=>	57286,
		8819	=>	57288,
		8820	=>	57290,
		8821	=>	57292,
		8822	=>	57294,
		8823	=>	57296,
		8824	=>	57298,
		8825	=>	57300,
		8826	=>	57302,
		8827	=>	57304,
		8828	=>	57307,
		8829	=>	57309,
		8830	=>	57311,
		8831	=>	57313,
		8832	=>	57315,
		8833	=>	57317,
		8834	=>	57319,
		8835	=>	57321,
		8836	=>	57323,
		8837	=>	57325,
		8838	=>	57327,
		8839	=>	57329,
		8840	=>	57331,
		8841	=>	57334,
		8842	=>	57336,
		8843	=>	57338,
		8844	=>	57340,
		8845	=>	57342,
		8846	=>	57344,
		8847	=>	57346,
		8848	=>	57348,
		8849	=>	57350,
		8850	=>	57352,
		8851	=>	57354,
		8852	=>	57356,
		8853	=>	57358,
		8854	=>	57361,
		8855	=>	57363,
		8856	=>	57365,
		8857	=>	57367,
		8858	=>	57369,
		8859	=>	57371,
		8860	=>	57373,
		8861	=>	57375,
		8862	=>	57377,
		8863	=>	57379,
		8864	=>	57381,
		8865	=>	57383,
		8866	=>	57385,
		8867	=>	57388,
		8868	=>	57390,
		8869	=>	57392,
		8870	=>	57394,
		8871	=>	57396,
		8872	=>	57398,
		8873	=>	57400,
		8874	=>	57402,
		8875	=>	57404,
		8876	=>	57406,
		8877	=>	57408,
		8878	=>	57410,
		8879	=>	57412,
		8880	=>	57414,
		8881	=>	57417,
		8882	=>	57419,
		8883	=>	57421,
		8884	=>	57423,
		8885	=>	57425,
		8886	=>	57427,
		8887	=>	57429,
		8888	=>	57431,
		8889	=>	57433,
		8890	=>	57435,
		8891	=>	57437,
		8892	=>	57439,
		8893	=>	57441,
		8894	=>	57443,
		8895	=>	57445,
		8896	=>	57448,
		8897	=>	57450,
		8898	=>	57452,
		8899	=>	57454,
		8900	=>	57456,
		8901	=>	57458,
		8902	=>	57460,
		8903	=>	57462,
		8904	=>	57464,
		8905	=>	57466,
		8906	=>	57468,
		8907	=>	57470,
		8908	=>	57472,
		8909	=>	57474,
		8910	=>	57476,
		8911	=>	57479,
		8912	=>	57481,
		8913	=>	57483,
		8914	=>	57485,
		8915	=>	57487,
		8916	=>	57489,
		8917	=>	57491,
		8918	=>	57493,
		8919	=>	57495,
		8920	=>	57497,
		8921	=>	57499,
		8922	=>	57501,
		8923	=>	57503,
		8924	=>	57505,
		8925	=>	57507,
		8926	=>	57509,
		8927	=>	57512,
		8928	=>	57514,
		8929	=>	57516,
		8930	=>	57518,
		8931	=>	57520,
		8932	=>	57522,
		8933	=>	57524,
		8934	=>	57526,
		8935	=>	57528,
		8936	=>	57530,
		8937	=>	57532,
		8938	=>	57534,
		8939	=>	57536,
		8940	=>	57538,
		8941	=>	57540,
		8942	=>	57542,
		8943	=>	57544,
		8944	=>	57546,
		8945	=>	57549,
		8946	=>	57551,
		8947	=>	57553,
		8948	=>	57555,
		8949	=>	57557,
		8950	=>	57559,
		8951	=>	57561,
		8952	=>	57563,
		8953	=>	57565,
		8954	=>	57567,
		8955	=>	57569,
		8956	=>	57571,
		8957	=>	57573,
		8958	=>	57575,
		8959	=>	57577,
		8960	=>	57579,
		8961	=>	57581,
		8962	=>	57583,
		8963	=>	57585,
		8964	=>	57588,
		8965	=>	57590,
		8966	=>	57592,
		8967	=>	57594,
		8968	=>	57596,
		8969	=>	57598,
		8970	=>	57600,
		8971	=>	57602,
		8972	=>	57604,
		8973	=>	57606,
		8974	=>	57608,
		8975	=>	57610,
		8976	=>	57612,
		8977	=>	57614,
		8978	=>	57616,
		8979	=>	57618,
		8980	=>	57620,
		8981	=>	57622,
		8982	=>	57624,
		8983	=>	57626,
		8984	=>	57629,
		8985	=>	57631,
		8986	=>	57633,
		8987	=>	57635,
		8988	=>	57637,
		8989	=>	57639,
		8990	=>	57641,
		8991	=>	57643,
		8992	=>	57645,
		8993	=>	57647,
		8994	=>	57649,
		8995	=>	57651,
		8996	=>	57653,
		8997	=>	57655,
		8998	=>	57657,
		8999	=>	57659,
		9000	=>	57661,
		9001	=>	57663,
		9002	=>	57665,
		9003	=>	57667,
		9004	=>	57669,
		9005	=>	57671,
		9006	=>	57673,
		9007	=>	57676,
		9008	=>	57678,
		9009	=>	57680,
		9010	=>	57682,
		9011	=>	57684,
		9012	=>	57686,
		9013	=>	57688,
		9014	=>	57690,
		9015	=>	57692,
		9016	=>	57694,
		9017	=>	57696,
		9018	=>	57698,
		9019	=>	57700,
		9020	=>	57702,
		9021	=>	57704,
		9022	=>	57706,
		9023	=>	57708,
		9024	=>	57710,
		9025	=>	57712,
		9026	=>	57714,
		9027	=>	57716,
		9028	=>	57718,
		9029	=>	57720,
		9030	=>	57722,
		9031	=>	57724,
		9032	=>	57726,
		9033	=>	57729,
		9034	=>	57731,
		9035	=>	57733,
		9036	=>	57735,
		9037	=>	57737,
		9038	=>	57739,
		9039	=>	57741,
		9040	=>	57743,
		9041	=>	57745,
		9042	=>	57747,
		9043	=>	57749,
		9044	=>	57751,
		9045	=>	57753,
		9046	=>	57755,
		9047	=>	57757,
		9048	=>	57759,
		9049	=>	57761,
		9050	=>	57763,
		9051	=>	57765,
		9052	=>	57767,
		9053	=>	57769,
		9054	=>	57771,
		9055	=>	57773,
		9056	=>	57775,
		9057	=>	57777,
		9058	=>	57779,
		9059	=>	57781,
		9060	=>	57783,
		9061	=>	57785,
		9062	=>	57787,
		9063	=>	57789,
		9064	=>	57792,
		9065	=>	57794,
		9066	=>	57796,
		9067	=>	57798,
		9068	=>	57800,
		9069	=>	57802,
		9070	=>	57804,
		9071	=>	57806,
		9072	=>	57808,
		9073	=>	57810,
		9074	=>	57812,
		9075	=>	57814,
		9076	=>	57816,
		9077	=>	57818,
		9078	=>	57820,
		9079	=>	57822,
		9080	=>	57824,
		9081	=>	57826,
		9082	=>	57828,
		9083	=>	57830,
		9084	=>	57832,
		9085	=>	57834,
		9086	=>	57836,
		9087	=>	57838,
		9088	=>	57840,
		9089	=>	57842,
		9090	=>	57844,
		9091	=>	57846,
		9092	=>	57848,
		9093	=>	57850,
		9094	=>	57852,
		9095	=>	57854,
		9096	=>	57856,
		9097	=>	57858,
		9098	=>	57860,
		9099	=>	57862,
		9100	=>	57864,
		9101	=>	57866,
		9102	=>	57868,
		9103	=>	57870,
		9104	=>	57872,
		9105	=>	57874,
		9106	=>	57876,
		9107	=>	57879,
		9108	=>	57881,
		9109	=>	57883,
		9110	=>	57885,
		9111	=>	57887,
		9112	=>	57889,
		9113	=>	57891,
		9114	=>	57893,
		9115	=>	57895,
		9116	=>	57897,
		9117	=>	57899,
		9118	=>	57901,
		9119	=>	57903,
		9120	=>	57905,
		9121	=>	57907,
		9122	=>	57909,
		9123	=>	57911,
		9124	=>	57913,
		9125	=>	57915,
		9126	=>	57917,
		9127	=>	57919,
		9128	=>	57921,
		9129	=>	57923,
		9130	=>	57925,
		9131	=>	57927,
		9132	=>	57929,
		9133	=>	57931,
		9134	=>	57933,
		9135	=>	57935,
		9136	=>	57937,
		9137	=>	57939,
		9138	=>	57941,
		9139	=>	57943,
		9140	=>	57945,
		9141	=>	57947,
		9142	=>	57949,
		9143	=>	57951,
		9144	=>	57953,
		9145	=>	57955,
		9146	=>	57957,
		9147	=>	57959,
		9148	=>	57961,
		9149	=>	57963,
		9150	=>	57965,
		9151	=>	57967,
		9152	=>	57969,
		9153	=>	57971,
		9154	=>	57973,
		9155	=>	57975,
		9156	=>	57977,
		9157	=>	57979,
		9158	=>	57981,
		9159	=>	57983,
		9160	=>	57985,
		9161	=>	57987,
		9162	=>	57989,
		9163	=>	57991,
		9164	=>	57993,
		9165	=>	57995,
		9166	=>	57997,
		9167	=>	57999,
		9168	=>	58001,
		9169	=>	58003,
		9170	=>	58005,
		9171	=>	58007,
		9172	=>	58009,
		9173	=>	58011,
		9174	=>	58013,
		9175	=>	58015,
		9176	=>	58017,
		9177	=>	58019,
		9178	=>	58021,
		9179	=>	58023,
		9180	=>	58025,
		9181	=>	58027,
		9182	=>	58029,
		9183	=>	58031,
		9184	=>	58033,
		9185	=>	58035,
		9186	=>	58037,
		9187	=>	58039,
		9188	=>	58041,
		9189	=>	58043,
		9190	=>	58045,
		9191	=>	58047,
		9192	=>	58049,
		9193	=>	58051,
		9194	=>	58053,
		9195	=>	58055,
		9196	=>	58057,
		9197	=>	58059,
		9198	=>	58061,
		9199	=>	58063,
		9200	=>	58065,
		9201	=>	58067,
		9202	=>	58069,
		9203	=>	58071,
		9204	=>	58073,
		9205	=>	58075,
		9206	=>	58077,
		9207	=>	58079,
		9208	=>	58081,
		9209	=>	58083,
		9210	=>	58085,
		9211	=>	58087,
		9212	=>	58089,
		9213	=>	58091,
		9214	=>	58093,
		9215	=>	58095,
		9216	=>	58097,
		9217	=>	58099,
		9218	=>	58101,
		9219	=>	58103,
		9220	=>	58105,
		9221	=>	58107,
		9222	=>	58109,
		9223	=>	58111,
		9224	=>	58113,
		9225	=>	58115,
		9226	=>	58117,
		9227	=>	58119,
		9228	=>	58121,
		9229	=>	58123,
		9230	=>	58125,
		9231	=>	58127,
		9232	=>	58129,
		9233	=>	58131,
		9234	=>	58133,
		9235	=>	58135,
		9236	=>	58137,
		9237	=>	58139,
		9238	=>	58141,
		9239	=>	58143,
		9240	=>	58145,
		9241	=>	58147,
		9242	=>	58149,
		9243	=>	58151,
		9244	=>	58153,
		9245	=>	58155,
		9246	=>	58157,
		9247	=>	58159,
		9248	=>	58161,
		9249	=>	58163,
		9250	=>	58165,
		9251	=>	58167,
		9252	=>	58169,
		9253	=>	58171,
		9254	=>	58173,
		9255	=>	58175,
		9256	=>	58177,
		9257	=>	58179,
		9258	=>	58181,
		9259	=>	58183,
		9260	=>	58185,
		9261	=>	58187,
		9262	=>	58189,
		9263	=>	58191,
		9264	=>	58193,
		9265	=>	58194,
		9266	=>	58196,
		9267	=>	58198,
		9268	=>	58200,
		9269	=>	58202,
		9270	=>	58204,
		9271	=>	58206,
		9272	=>	58208,
		9273	=>	58210,
		9274	=>	58212,
		9275	=>	58214,
		9276	=>	58216,
		9277	=>	58218,
		9278	=>	58220,
		9279	=>	58222,
		9280	=>	58224,
		9281	=>	58226,
		9282	=>	58228,
		9283	=>	58230,
		9284	=>	58232,
		9285	=>	58234,
		9286	=>	58236,
		9287	=>	58238,
		9288	=>	58240,
		9289	=>	58242,
		9290	=>	58244,
		9291	=>	58246,
		9292	=>	58248,
		9293	=>	58250,
		9294	=>	58252,
		9295	=>	58254,
		9296	=>	58256,
		9297	=>	58258,
		9298	=>	58260,
		9299	=>	58262,
		9300	=>	58264,
		9301	=>	58266,
		9302	=>	58268,
		9303	=>	58270,
		9304	=>	58272,
		9305	=>	58274,
		9306	=>	58276,
		9307	=>	58278,
		9308	=>	58279,
		9309	=>	58281,
		9310	=>	58283,
		9311	=>	58285,
		9312	=>	58287,
		9313	=>	58289,
		9314	=>	58291,
		9315	=>	58293,
		9316	=>	58295,
		9317	=>	58297,
		9318	=>	58299,
		9319	=>	58301,
		9320	=>	58303,
		9321	=>	58305,
		9322	=>	58307,
		9323	=>	58309,
		9324	=>	58311,
		9325	=>	58313,
		9326	=>	58315,
		9327	=>	58317,
		9328	=>	58319,
		9329	=>	58321,
		9330	=>	58323,
		9331	=>	58325,
		9332	=>	58327,
		9333	=>	58329,
		9334	=>	58331,
		9335	=>	58333,
		9336	=>	58335,
		9337	=>	58337,
		9338	=>	58339,
		9339	=>	58340,
		9340	=>	58342,
		9341	=>	58344,
		9342	=>	58346,
		9343	=>	58348,
		9344	=>	58350,
		9345	=>	58352,
		9346	=>	58354,
		9347	=>	58356,
		9348	=>	58358,
		9349	=>	58360,
		9350	=>	58362,
		9351	=>	58364,
		9352	=>	58366,
		9353	=>	58368,
		9354	=>	58370,
		9355	=>	58372,
		9356	=>	58374,
		9357	=>	58376,
		9358	=>	58378,
		9359	=>	58380,
		9360	=>	58382,
		9361	=>	58384,
		9362	=>	58386,
		9363	=>	58388,
		9364	=>	58390,
		9365	=>	58391,
		9366	=>	58393,
		9367	=>	58395,
		9368	=>	58397,
		9369	=>	58399,
		9370	=>	58401,
		9371	=>	58403,
		9372	=>	58405,
		9373	=>	58407,
		9374	=>	58409,
		9375	=>	58411,
		9376	=>	58413,
		9377	=>	58415,
		9378	=>	58417,
		9379	=>	58419,
		9380	=>	58421,
		9381	=>	58423,
		9382	=>	58425,
		9383	=>	58427,
		9384	=>	58429,
		9385	=>	58431,
		9386	=>	58433,
		9387	=>	58434,
		9388	=>	58436,
		9389	=>	58438,
		9390	=>	58440,
		9391	=>	58442,
		9392	=>	58444,
		9393	=>	58446,
		9394	=>	58448,
		9395	=>	58450,
		9396	=>	58452,
		9397	=>	58454,
		9398	=>	58456,
		9399	=>	58458,
		9400	=>	58460,
		9401	=>	58462,
		9402	=>	58464,
		9403	=>	58466,
		9404	=>	58468,
		9405	=>	58470,
		9406	=>	58472,
		9407	=>	58474,
		9408	=>	58475,
		9409	=>	58477,
		9410	=>	58479,
		9411	=>	58481,
		9412	=>	58483,
		9413	=>	58485,
		9414	=>	58487,
		9415	=>	58489,
		9416	=>	58491,
		9417	=>	58493,
		9418	=>	58495,
		9419	=>	58497,
		9420	=>	58499,
		9421	=>	58501,
		9422	=>	58503,
		9423	=>	58505,
		9424	=>	58507,
		9425	=>	58509,
		9426	=>	58510,
		9427	=>	58512,
		9428	=>	58514,
		9429	=>	58516,
		9430	=>	58518,
		9431	=>	58520,
		9432	=>	58522,
		9433	=>	58524,
		9434	=>	58526,
		9435	=>	58528,
		9436	=>	58530,
		9437	=>	58532,
		9438	=>	58534,
		9439	=>	58536,
		9440	=>	58538,
		9441	=>	58540,
		9442	=>	58542,
		9443	=>	58543,
		9444	=>	58545,
		9445	=>	58547,
		9446	=>	58549,
		9447	=>	58551,
		9448	=>	58553,
		9449	=>	58555,
		9450	=>	58557,
		9451	=>	58559,
		9452	=>	58561,
		9453	=>	58563,
		9454	=>	58565,
		9455	=>	58567,
		9456	=>	58569,
		9457	=>	58571,
		9458	=>	58573,
		9459	=>	58574,
		9460	=>	58576,
		9461	=>	58578,
		9462	=>	58580,
		9463	=>	58582,
		9464	=>	58584,
		9465	=>	58586,
		9466	=>	58588,
		9467	=>	58590,
		9468	=>	58592,
		9469	=>	58594,
		9470	=>	58596,
		9471	=>	58598,
		9472	=>	58600,
		9473	=>	58602,
		9474	=>	58604,
		9475	=>	58605,
		9476	=>	58607,
		9477	=>	58609,
		9478	=>	58611,
		9479	=>	58613,
		9480	=>	58615,
		9481	=>	58617,
		9482	=>	58619,
		9483	=>	58621,
		9484	=>	58623,
		9485	=>	58625,
		9486	=>	58627,
		9487	=>	58629,
		9488	=>	58631,
		9489	=>	58632,
		9490	=>	58634,
		9491	=>	58636,
		9492	=>	58638,
		9493	=>	58640,
		9494	=>	58642,
		9495	=>	58644,
		9496	=>	58646,
		9497	=>	58648,
		9498	=>	58650,
		9499	=>	58652,
		9500	=>	58654,
		9501	=>	58656,
		9502	=>	58658,
		9503	=>	58659,
		9504	=>	58661,
		9505	=>	58663,
		9506	=>	58665,
		9507	=>	58667,
		9508	=>	58669,
		9509	=>	58671,
		9510	=>	58673,
		9511	=>	58675,
		9512	=>	58677,
		9513	=>	58679,
		9514	=>	58681,
		9515	=>	58683,
		9516	=>	58684,
		9517	=>	58686,
		9518	=>	58688,
		9519	=>	58690,
		9520	=>	58692,
		9521	=>	58694,
		9522	=>	58696,
		9523	=>	58698,
		9524	=>	58700,
		9525	=>	58702,
		9526	=>	58704,
		9527	=>	58706,
		9528	=>	58708,
		9529	=>	58709,
		9530	=>	58711,
		9531	=>	58713,
		9532	=>	58715,
		9533	=>	58717,
		9534	=>	58719,
		9535	=>	58721,
		9536	=>	58723,
		9537	=>	58725,
		9538	=>	58727,
		9539	=>	58729,
		9540	=>	58731,
		9541	=>	58732,
		9542	=>	58734,
		9543	=>	58736,
		9544	=>	58738,
		9545	=>	58740,
		9546	=>	58742,
		9547	=>	58744,
		9548	=>	58746,
		9549	=>	58748,
		9550	=>	58750,
		9551	=>	58752,
		9552	=>	58754,
		9553	=>	58755,
		9554	=>	58757,
		9555	=>	58759,
		9556	=>	58761,
		9557	=>	58763,
		9558	=>	58765,
		9559	=>	58767,
		9560	=>	58769,
		9561	=>	58771,
		9562	=>	58773,
		9563	=>	58775,
		9564	=>	58776,
		9565	=>	58778,
		9566	=>	58780,
		9567	=>	58782,
		9568	=>	58784,
		9569	=>	58786,
		9570	=>	58788,
		9571	=>	58790,
		9572	=>	58792,
		9573	=>	58794,
		9574	=>	58796,
		9575	=>	58797,
		9576	=>	58799,
		9577	=>	58801,
		9578	=>	58803,
		9579	=>	58805,
		9580	=>	58807,
		9581	=>	58809,
		9582	=>	58811,
		9583	=>	58813,
		9584	=>	58815,
		9585	=>	58817,
		9586	=>	58818,
		9587	=>	58820,
		9588	=>	58822,
		9589	=>	58824,
		9590	=>	58826,
		9591	=>	58828,
		9592	=>	58830,
		9593	=>	58832,
		9594	=>	58834,
		9595	=>	58836,
		9596	=>	58837,
		9597	=>	58839,
		9598	=>	58841,
		9599	=>	58843,
		9600	=>	58845,
		9601	=>	58847,
		9602	=>	58849,
		9603	=>	58851,
		9604	=>	58853,
		9605	=>	58855,
		9606	=>	58856,
		9607	=>	58858,
		9608	=>	58860,
		9609	=>	58862,
		9610	=>	58864,
		9611	=>	58866,
		9612	=>	58868,
		9613	=>	58870,
		9614	=>	58872,
		9615	=>	58874,
		9616	=>	58875,
		9617	=>	58877,
		9618	=>	58879,
		9619	=>	58881,
		9620	=>	58883,
		9621	=>	58885,
		9622	=>	58887,
		9623	=>	58889,
		9624	=>	58891,
		9625	=>	58893,
		9626	=>	58894,
		9627	=>	58896,
		9628	=>	58898,
		9629	=>	58900,
		9630	=>	58902,
		9631	=>	58904,
		9632	=>	58906,
		9633	=>	58908,
		9634	=>	58910,
		9635	=>	58912,
		9636	=>	58913,
		9637	=>	58915,
		9638	=>	58917,
		9639	=>	58919,
		9640	=>	58921,
		9641	=>	58923,
		9642	=>	58925,
		9643	=>	58927,
		9644	=>	58929,
		9645	=>	58930,
		9646	=>	58932,
		9647	=>	58934,
		9648	=>	58936,
		9649	=>	58938,
		9650	=>	58940,
		9651	=>	58942,
		9652	=>	58944,
		9653	=>	58946,
		9654	=>	58947,
		9655	=>	58949,
		9656	=>	58951,
		9657	=>	58953,
		9658	=>	58955,
		9659	=>	58957,
		9660	=>	58959,
		9661	=>	58961,
		9662	=>	58963,
		9663	=>	58964,
		9664	=>	58966,
		9665	=>	58968,
		9666	=>	58970,
		9667	=>	58972,
		9668	=>	58974,
		9669	=>	58976,
		9670	=>	58978,
		9671	=>	58980,
		9672	=>	58981,
		9673	=>	58983,
		9674	=>	58985,
		9675	=>	58987,
		9676	=>	58989,
		9677	=>	58991,
		9678	=>	58993,
		9679	=>	58995,
		9680	=>	58996,
		9681	=>	58998,
		9682	=>	59000,
		9683	=>	59002,
		9684	=>	59004,
		9685	=>	59006,
		9686	=>	59008,
		9687	=>	59010,
		9688	=>	59012,
		9689	=>	59013,
		9690	=>	59015,
		9691	=>	59017,
		9692	=>	59019,
		9693	=>	59021,
		9694	=>	59023,
		9695	=>	59025,
		9696	=>	59027,
		9697	=>	59028,
		9698	=>	59030,
		9699	=>	59032,
		9700	=>	59034,
		9701	=>	59036,
		9702	=>	59038,
		9703	=>	59040,
		9704	=>	59042,
		9705	=>	59043,
		9706	=>	59045,
		9707	=>	59047,
		9708	=>	59049,
		9709	=>	59051,
		9710	=>	59053,
		9711	=>	59055,
		9712	=>	59057,
		9713	=>	59059,
		9714	=>	59060,
		9715	=>	59062,
		9716	=>	59064,
		9717	=>	59066,
		9718	=>	59068,
		9719	=>	59070,
		9720	=>	59072,
		9721	=>	59073,
		9722	=>	59075,
		9723	=>	59077,
		9724	=>	59079,
		9725	=>	59081,
		9726	=>	59083,
		9727	=>	59085,
		9728	=>	59087,
		9729	=>	59088,
		9730	=>	59090,
		9731	=>	59092,
		9732	=>	59094,
		9733	=>	59096,
		9734	=>	59098,
		9735	=>	59100,
		9736	=>	59102,
		9737	=>	59103,
		9738	=>	59105,
		9739	=>	59107,
		9740	=>	59109,
		9741	=>	59111,
		9742	=>	59113,
		9743	=>	59115,
		9744	=>	59117,
		9745	=>	59118,
		9746	=>	59120,
		9747	=>	59122,
		9748	=>	59124,
		9749	=>	59126,
		9750	=>	59128,
		9751	=>	59130,
		9752	=>	59131,
		9753	=>	59133,
		9754	=>	59135,
		9755	=>	59137,
		9756	=>	59139,
		9757	=>	59141,
		9758	=>	59143,
		9759	=>	59145,
		9760	=>	59146,
		9761	=>	59148,
		9762	=>	59150,
		9763	=>	59152,
		9764	=>	59154,
		9765	=>	59156,
		9766	=>	59158,
		9767	=>	59159,
		9768	=>	59161,
		9769	=>	59163,
		9770	=>	59165,
		9771	=>	59167,
		9772	=>	59169,
		9773	=>	59171,
		9774	=>	59172,
		9775	=>	59174,
		9776	=>	59176,
		9777	=>	59178,
		9778	=>	59180,
		9779	=>	59182,
		9780	=>	59184,
		9781	=>	59185,
		9782	=>	59187,
		9783	=>	59189,
		9784	=>	59191,
		9785	=>	59193,
		9786	=>	59195,
		9787	=>	59197,
		9788	=>	59198,
		9789	=>	59200,
		9790	=>	59202,
		9791	=>	59204,
		9792	=>	59206,
		9793	=>	59208,
		9794	=>	59210,
		9795	=>	59211,
		9796	=>	59213,
		9797	=>	59215,
		9798	=>	59217,
		9799	=>	59219,
		9800	=>	59221,
		9801	=>	59223,
		9802	=>	59224,
		9803	=>	59226,
		9804	=>	59228,
		9805	=>	59230,
		9806	=>	59232,
		9807	=>	59234,
		9808	=>	59236,
		9809	=>	59237,
		9810	=>	59239,
		9811	=>	59241,
		9812	=>	59243,
		9813	=>	59245,
		9814	=>	59247,
		9815	=>	59248,
		9816	=>	59250,
		9817	=>	59252,
		9818	=>	59254,
		9819	=>	59256,
		9820	=>	59258,
		9821	=>	59260,
		9822	=>	59261,
		9823	=>	59263,
		9824	=>	59265,
		9825	=>	59267,
		9826	=>	59269,
		9827	=>	59271,
		9828	=>	59273,
		9829	=>	59274,
		9830	=>	59276,
		9831	=>	59278,
		9832	=>	59280,
		9833	=>	59282,
		9834	=>	59284,
		9835	=>	59285,
		9836	=>	59287,
		9837	=>	59289,
		9838	=>	59291,
		9839	=>	59293,
		9840	=>	59295,
		9841	=>	59297,
		9842	=>	59298,
		9843	=>	59300,
		9844	=>	59302,
		9845	=>	59304,
		9846	=>	59306,
		9847	=>	59308,
		9848	=>	59309,
		9849	=>	59311,
		9850	=>	59313,
		9851	=>	59315,
		9852	=>	59317,
		9853	=>	59319,
		9854	=>	59320,
		9855	=>	59322,
		9856	=>	59324,
		9857	=>	59326,
		9858	=>	59328,
		9859	=>	59330,
		9860	=>	59332,
		9861	=>	59333,
		9862	=>	59335,
		9863	=>	59337,
		9864	=>	59339,
		9865	=>	59341,
		9866	=>	59343,
		9867	=>	59344,
		9868	=>	59346,
		9869	=>	59348,
		9870	=>	59350,
		9871	=>	59352,
		9872	=>	59354,
		9873	=>	59355,
		9874	=>	59357,
		9875	=>	59359,
		9876	=>	59361,
		9877	=>	59363,
		9878	=>	59365,
		9879	=>	59366,
		9880	=>	59368,
		9881	=>	59370,
		9882	=>	59372,
		9883	=>	59374,
		9884	=>	59376,
		9885	=>	59377,
		9886	=>	59379,
		9887	=>	59381,
		9888	=>	59383,
		9889	=>	59385,
		9890	=>	59387,
		9891	=>	59388,
		9892	=>	59390,
		9893	=>	59392,
		9894	=>	59394,
		9895	=>	59396,
		9896	=>	59398,
		9897	=>	59399,
		9898	=>	59401,
		9899	=>	59403,
		9900	=>	59405,
		9901	=>	59407,
		9902	=>	59409,
		9903	=>	59410,
		9904	=>	59412,
		9905	=>	59414,
		9906	=>	59416,
		9907	=>	59418,
		9908	=>	59420,
		9909	=>	59421,
		9910	=>	59423,
		9911	=>	59425,
		9912	=>	59427,
		9913	=>	59429,
		9914	=>	59430,
		9915	=>	59432,
		9916	=>	59434,
		9917	=>	59436,
		9918	=>	59438,
		9919	=>	59440,
		9920	=>	59441,
		9921	=>	59443,
		9922	=>	59445,
		9923	=>	59447,
		9924	=>	59449,
		9925	=>	59451,
		9926	=>	59452,
		9927	=>	59454,
		9928	=>	59456,
		9929	=>	59458,
		9930	=>	59460,
		9931	=>	59461,
		9932	=>	59463,
		9933	=>	59465,
		9934	=>	59467,
		9935	=>	59469,
		9936	=>	59471,
		9937	=>	59472,
		9938	=>	59474,
		9939	=>	59476,
		9940	=>	59478,
		9941	=>	59480,
		9942	=>	59482,
		9943	=>	59483,
		9944	=>	59485,
		9945	=>	59487,
		9946	=>	59489,
		9947	=>	59491,
		9948	=>	59492,
		9949	=>	59494,
		9950	=>	59496,
		9951	=>	59498,
		9952	=>	59500,
		9953	=>	59502,
		9954	=>	59503,
		9955	=>	59505,
		9956	=>	59507,
		9957	=>	59509,
		9958	=>	59511,
		9959	=>	59512,
		9960	=>	59514,
		9961	=>	59516,
		9962	=>	59518,
		9963	=>	59520,
		9964	=>	59521,
		9965	=>	59523,
		9966	=>	59525,
		9967	=>	59527,
		9968	=>	59529,
		9969	=>	59531,
		9970	=>	59532,
		9971	=>	59534,
		9972	=>	59536,
		9973	=>	59538,
		9974	=>	59540,
		9975	=>	59541,
		9976	=>	59543,
		9977	=>	59545,
		9978	=>	59547,
		9979	=>	59549,
		9980	=>	59550,
		9981	=>	59552,
		9982	=>	59554,
		9983	=>	59556,
		9984	=>	59558,
		9985	=>	59560,
		9986	=>	59561,
		9987	=>	59563,
		9988	=>	59565,
		9989	=>	59567,
		9990	=>	59569,
		9991	=>	59570,
		9992	=>	59572,
		9993	=>	59574,
		9994	=>	59576,
		9995	=>	59578,
		9996	=>	59579,
		9997	=>	59581,
		9998	=>	59583,
		9999	=>	59585,
		10000	=>	59587,
		10001	=>	59588,
		10002	=>	59590,
		10003	=>	59592,
		10004	=>	59594,
		10005	=>	59596,
		10006	=>	59597,
		10007	=>	59599,
		10008	=>	59601,
		10009	=>	59603,
		10010	=>	59605,
		10011	=>	59606,
		10012	=>	59608,
		10013	=>	59610,
		10014	=>	59612,
		10015	=>	59614,
		10016	=>	59615,
		10017	=>	59617,
		10018	=>	59619,
		10019	=>	59621,
		10020	=>	59623,
		10021	=>	59624,
		10022	=>	59626,
		10023	=>	59628,
		10024	=>	59630,
		10025	=>	59632,
		10026	=>	59633,
		10027	=>	59635,
		10028	=>	59637,
		10029	=>	59639,
		10030	=>	59641,
		10031	=>	59642,
		10032	=>	59644,
		10033	=>	59646,
		10034	=>	59648,
		10035	=>	59650,
		10036	=>	59651,
		10037	=>	59653,
		10038	=>	59655,
		10039	=>	59657,
		10040	=>	59659,
		10041	=>	59660,
		10042	=>	59662,
		10043	=>	59664,
		10044	=>	59666,
		10045	=>	59668,
		10046	=>	59669,
		10047	=>	59671,
		10048	=>	59673,
		10049	=>	59675,
		10050	=>	59677,
		10051	=>	59678,
		10052	=>	59680,
		10053	=>	59682,
		10054	=>	59684,
		10055	=>	59686,
		10056	=>	59687,
		10057	=>	59689,
		10058	=>	59691,
		10059	=>	59693,
		10060	=>	59694,
		10061	=>	59696,
		10062	=>	59698,
		10063	=>	59700,
		10064	=>	59702,
		10065	=>	59703,
		10066	=>	59705,
		10067	=>	59707,
		10068	=>	59709,
		10069	=>	59711,
		10070	=>	59712,
		10071	=>	59714,
		10072	=>	59716,
		10073	=>	59718,
		10074	=>	59720,
		10075	=>	59721,
		10076	=>	59723,
		10077	=>	59725,
		10078	=>	59727,
		10079	=>	59728,
		10080	=>	59730,
		10081	=>	59732,
		10082	=>	59734,
		10083	=>	59736,
		10084	=>	59737,
		10085	=>	59739,
		10086	=>	59741,
		10087	=>	59743,
		10088	=>	59745,
		10089	=>	59746,
		10090	=>	59748,
		10091	=>	59750,
		10092	=>	59752,
		10093	=>	59753,
		10094	=>	59755,
		10095	=>	59757,
		10096	=>	59759,
		10097	=>	59761,
		10098	=>	59762,
		10099	=>	59764,
		10100	=>	59766,
		10101	=>	59768,
		10102	=>	59769,
		10103	=>	59771,
		10104	=>	59773,
		10105	=>	59775,
		10106	=>	59777,
		10107	=>	59778,
		10108	=>	59780,
		10109	=>	59782,
		10110	=>	59784,
		10111	=>	59785,
		10112	=>	59787,
		10113	=>	59789,
		10114	=>	59791,
		10115	=>	59793,
		10116	=>	59794,
		10117	=>	59796,
		10118	=>	59798,
		10119	=>	59800,
		10120	=>	59801,
		10121	=>	59803,
		10122	=>	59805,
		10123	=>	59807,
		10124	=>	59809,
		10125	=>	59810,
		10126	=>	59812,
		10127	=>	59814,
		10128	=>	59816,
		10129	=>	59817,
		10130	=>	59819,
		10131	=>	59821,
		10132	=>	59823,
		10133	=>	59824,
		10134	=>	59826,
		10135	=>	59828,
		10136	=>	59830,
		10137	=>	59832,
		10138	=>	59833,
		10139	=>	59835,
		10140	=>	59837,
		10141	=>	59839,
		10142	=>	59840,
		10143	=>	59842,
		10144	=>	59844,
		10145	=>	59846,
		10146	=>	59848,
		10147	=>	59849,
		10148	=>	59851,
		10149	=>	59853,
		10150	=>	59855,
		10151	=>	59856,
		10152	=>	59858,
		10153	=>	59860,
		10154	=>	59862,
		10155	=>	59863,
		10156	=>	59865,
		10157	=>	59867,
		10158	=>	59869,
		10159	=>	59870,
		10160	=>	59872,
		10161	=>	59874,
		10162	=>	59876,
		10163	=>	59878,
		10164	=>	59879,
		10165	=>	59881,
		10166	=>	59883,
		10167	=>	59885,
		10168	=>	59886,
		10169	=>	59888,
		10170	=>	59890,
		10171	=>	59892,
		10172	=>	59893,
		10173	=>	59895,
		10174	=>	59897,
		10175	=>	59899,
		10176	=>	59900,
		10177	=>	59902,
		10178	=>	59904,
		10179	=>	59906,
		10180	=>	59908,
		10181	=>	59909,
		10182	=>	59911,
		10183	=>	59913,
		10184	=>	59915,
		10185	=>	59916,
		10186	=>	59918,
		10187	=>	59920,
		10188	=>	59922,
		10189	=>	59923,
		10190	=>	59925,
		10191	=>	59927,
		10192	=>	59929,
		10193	=>	59930,
		10194	=>	59932,
		10195	=>	59934,
		10196	=>	59936,
		10197	=>	59937,
		10198	=>	59939,
		10199	=>	59941,
		10200	=>	59943,
		10201	=>	59944,
		10202	=>	59946,
		10203	=>	59948,
		10204	=>	59950,
		10205	=>	59951,
		10206	=>	59953,
		10207	=>	59955,
		10208	=>	59957,
		10209	=>	59958,
		10210	=>	59960,
		10211	=>	59962,
		10212	=>	59964,
		10213	=>	59965,
		10214	=>	59967,
		10215	=>	59969,
		10216	=>	59971,
		10217	=>	59972,
		10218	=>	59974,
		10219	=>	59976,
		10220	=>	59978,
		10221	=>	59979,
		10222	=>	59981,
		10223	=>	59983,
		10224	=>	59985,
		10225	=>	59986,
		10226	=>	59988,
		10227	=>	59990,
		10228	=>	59992,
		10229	=>	59993,
		10230	=>	59995,
		10231	=>	59997,
		10232	=>	59999,
		10233	=>	60000,
		10234	=>	60002,
		10235	=>	60004,
		10236	=>	60006,
		10237	=>	60007,
		10238	=>	60009,
		10239	=>	60011,
		10240	=>	60013,
		10241	=>	60014,
		10242	=>	60016,
		10243	=>	60018,
		10244	=>	60020,
		10245	=>	60021,
		10246	=>	60023,
		10247	=>	60025,
		10248	=>	60027,
		10249	=>	60028,
		10250	=>	60030,
		10251	=>	60032,
		10252	=>	60034,
		10253	=>	60035,
		10254	=>	60037,
		10255	=>	60039,
		10256	=>	60041,
		10257	=>	60042,
		10258	=>	60044,
		10259	=>	60046,
		10260	=>	60048,
		10261	=>	60049,
		10262	=>	60051,
		10263	=>	60053,
		10264	=>	60054,
		10265	=>	60056,
		10266	=>	60058,
		10267	=>	60060,
		10268	=>	60061,
		10269	=>	60063,
		10270	=>	60065,
		10271	=>	60067,
		10272	=>	60068,
		10273	=>	60070,
		10274	=>	60072,
		10275	=>	60074,
		10276	=>	60075,
		10277	=>	60077,
		10278	=>	60079,
		10279	=>	60081,
		10280	=>	60082,
		10281	=>	60084,
		10282	=>	60086,
		10283	=>	60087,
		10284	=>	60089,
		10285	=>	60091,
		10286	=>	60093,
		10287	=>	60094,
		10288	=>	60096,
		10289	=>	60098,
		10290	=>	60100,
		10291	=>	60101,
		10292	=>	60103,
		10293	=>	60105,
		10294	=>	60107,
		10295	=>	60108,
		10296	=>	60110,
		10297	=>	60112,
		10298	=>	60113,
		10299	=>	60115,
		10300	=>	60117,
		10301	=>	60119,
		10302	=>	60120,
		10303	=>	60122,
		10304	=>	60124,
		10305	=>	60126,
		10306	=>	60127,
		10307	=>	60129,
		10308	=>	60131,
		10309	=>	60133,
		10310	=>	60134,
		10311	=>	60136,
		10312	=>	60138,
		10313	=>	60139,
		10314	=>	60141,
		10315	=>	60143,
		10316	=>	60145,
		10317	=>	60146,
		10318	=>	60148,
		10319	=>	60150,
		10320	=>	60152,
		10321	=>	60153,
		10322	=>	60155,
		10323	=>	60157,
		10324	=>	60158,
		10325	=>	60160,
		10326	=>	60162,
		10327	=>	60164,
		10328	=>	60165,
		10329	=>	60167,
		10330	=>	60169,
		10331	=>	60170,
		10332	=>	60172,
		10333	=>	60174,
		10334	=>	60176,
		10335	=>	60177,
		10336	=>	60179,
		10337	=>	60181,
		10338	=>	60183,
		10339	=>	60184,
		10340	=>	60186,
		10341	=>	60188,
		10342	=>	60189,
		10343	=>	60191,
		10344	=>	60193,
		10345	=>	60195,
		10346	=>	60196,
		10347	=>	60198,
		10348	=>	60200,
		10349	=>	60201,
		10350	=>	60203,
		10351	=>	60205,
		10352	=>	60207,
		10353	=>	60208,
		10354	=>	60210,
		10355	=>	60212,
		10356	=>	60213,
		10357	=>	60215,
		10358	=>	60217,
		10359	=>	60219,
		10360	=>	60220,
		10361	=>	60222,
		10362	=>	60224,
		10363	=>	60225,
		10364	=>	60227,
		10365	=>	60229,
		10366	=>	60231,
		10367	=>	60232,
		10368	=>	60234,
		10369	=>	60236,
		10370	=>	60237,
		10371	=>	60239,
		10372	=>	60241,
		10373	=>	60243,
		10374	=>	60244,
		10375	=>	60246,
		10376	=>	60248,
		10377	=>	60249,
		10378	=>	60251,
		10379	=>	60253,
		10380	=>	60255,
		10381	=>	60256,
		10382	=>	60258,
		10383	=>	60260,
		10384	=>	60261,
		10385	=>	60263,
		10386	=>	60265,
		10387	=>	60267,
		10388	=>	60268,
		10389	=>	60270,
		10390	=>	60272,
		10391	=>	60273,
		10392	=>	60275,
		10393	=>	60277,
		10394	=>	60278,
		10395	=>	60280,
		10396	=>	60282,
		10397	=>	60284,
		10398	=>	60285,
		10399	=>	60287,
		10400	=>	60289,
		10401	=>	60290,
		10402	=>	60292,
		10403	=>	60294,
		10404	=>	60296,
		10405	=>	60297,
		10406	=>	60299,
		10407	=>	60301,
		10408	=>	60302,
		10409	=>	60304,
		10410	=>	60306,
		10411	=>	60307,
		10412	=>	60309,
		10413	=>	60311,
		10414	=>	60313,
		10415	=>	60314,
		10416	=>	60316,
		10417	=>	60318,
		10418	=>	60319,
		10419	=>	60321,
		10420	=>	60323,
		10421	=>	60324,
		10422	=>	60326,
		10423	=>	60328,
		10424	=>	60330,
		10425	=>	60331,
		10426	=>	60333,
		10427	=>	60335,
		10428	=>	60336,
		10429	=>	60338,
		10430	=>	60340,
		10431	=>	60341,
		10432	=>	60343,
		10433	=>	60345,
		10434	=>	60347,
		10435	=>	60348,
		10436	=>	60350,
		10437	=>	60352,
		10438	=>	60353,
		10439	=>	60355,
		10440	=>	60357,
		10441	=>	60358,
		10442	=>	60360,
		10443	=>	60362,
		10444	=>	60363,
		10445	=>	60365,
		10446	=>	60367,
		10447	=>	60369,
		10448	=>	60370,
		10449	=>	60372,
		10450	=>	60374,
		10451	=>	60375,
		10452	=>	60377,
		10453	=>	60379,
		10454	=>	60380,
		10455	=>	60382,
		10456	=>	60384,
		10457	=>	60385,
		10458	=>	60387,
		10459	=>	60389,
		10460	=>	60391,
		10461	=>	60392,
		10462	=>	60394,
		10463	=>	60396,
		10464	=>	60397,
		10465	=>	60399,
		10466	=>	60401,
		10467	=>	60402,
		10468	=>	60404,
		10469	=>	60406,
		10470	=>	60407,
		10471	=>	60409,
		10472	=>	60411,
		10473	=>	60413,
		10474	=>	60414,
		10475	=>	60416,
		10476	=>	60418,
		10477	=>	60419,
		10478	=>	60421,
		10479	=>	60423,
		10480	=>	60424,
		10481	=>	60426,
		10482	=>	60428,
		10483	=>	60429,
		10484	=>	60431,
		10485	=>	60433,
		10486	=>	60434,
		10487	=>	60436,
		10488	=>	60438,
		10489	=>	60439,
		10490	=>	60441,
		10491	=>	60443,
		10492	=>	60445,
		10493	=>	60446,
		10494	=>	60448,
		10495	=>	60450,
		10496	=>	60451,
		10497	=>	60453,
		10498	=>	60455,
		10499	=>	60456,
		10500	=>	60458,
		10501	=>	60460,
		10502	=>	60461,
		10503	=>	60463,
		10504	=>	60465,
		10505	=>	60466,
		10506	=>	60468,
		10507	=>	60470,
		10508	=>	60471,
		10509	=>	60473,
		10510	=>	60475,
		10511	=>	60476,
		10512	=>	60478,
		10513	=>	60480,
		10514	=>	60481,
		10515	=>	60483,
		10516	=>	60485,
		10517	=>	60486,
		10518	=>	60488,
		10519	=>	60490,
		10520	=>	60492,
		10521	=>	60493,
		10522	=>	60495,
		10523	=>	60497,
		10524	=>	60498,
		10525	=>	60500,
		10526	=>	60502,
		10527	=>	60503,
		10528	=>	60505,
		10529	=>	60507,
		10530	=>	60508,
		10531	=>	60510,
		10532	=>	60512,
		10533	=>	60513,
		10534	=>	60515,
		10535	=>	60517,
		10536	=>	60518,
		10537	=>	60520,
		10538	=>	60522,
		10539	=>	60523,
		10540	=>	60525,
		10541	=>	60527,
		10542	=>	60528,
		10543	=>	60530,
		10544	=>	60532,
		10545	=>	60533,
		10546	=>	60535,
		10547	=>	60537,
		10548	=>	60538,
		10549	=>	60540,
		10550	=>	60542,
		10551	=>	60543,
		10552	=>	60545,
		10553	=>	60547,
		10554	=>	60548,
		10555	=>	60550,
		10556	=>	60552,
		10557	=>	60553,
		10558	=>	60555,
		10559	=>	60557,
		10560	=>	60558,
		10561	=>	60560,
		10562	=>	60562,
		10563	=>	60563,
		10564	=>	60565,
		10565	=>	60567,
		10566	=>	60568,
		10567	=>	60570,
		10568	=>	60572,
		10569	=>	60573,
		10570	=>	60575,
		10571	=>	60577,
		10572	=>	60578,
		10573	=>	60580,
		10574	=>	60582,
		10575	=>	60583,
		10576	=>	60585,
		10577	=>	60587,
		10578	=>	60588,
		10579	=>	60590,
		10580	=>	60592,
		10581	=>	60593,
		10582	=>	60595,
		10583	=>	60596,
		10584	=>	60598,
		10585	=>	60600,
		10586	=>	60601,
		10587	=>	60603,
		10588	=>	60605,
		10589	=>	60606,
		10590	=>	60608,
		10591	=>	60610,
		10592	=>	60611,
		10593	=>	60613,
		10594	=>	60615,
		10595	=>	60616,
		10596	=>	60618,
		10597	=>	60620,
		10598	=>	60621,
		10599	=>	60623,
		10600	=>	60625,
		10601	=>	60626,
		10602	=>	60628,
		10603	=>	60630,
		10604	=>	60631,
		10605	=>	60633,
		10606	=>	60635,
		10607	=>	60636,
		10608	=>	60638,
		10609	=>	60640,
		10610	=>	60641,
		10611	=>	60643,
		10612	=>	60644,
		10613	=>	60646,
		10614	=>	60648,
		10615	=>	60649,
		10616	=>	60651,
		10617	=>	60653,
		10618	=>	60654,
		10619	=>	60656,
		10620	=>	60658,
		10621	=>	60659,
		10622	=>	60661,
		10623	=>	60663,
		10624	=>	60664,
		10625	=>	60666,
		10626	=>	60668,
		10627	=>	60669,
		10628	=>	60671,
		10629	=>	60673,
		10630	=>	60674,
		10631	=>	60676,
		10632	=>	60677,
		10633	=>	60679,
		10634	=>	60681,
		10635	=>	60682,
		10636	=>	60684,
		10637	=>	60686,
		10638	=>	60687,
		10639	=>	60689,
		10640	=>	60691,
		10641	=>	60692,
		10642	=>	60694,
		10643	=>	60696,
		10644	=>	60697,
		10645	=>	60699,
		10646	=>	60700,
		10647	=>	60702,
		10648	=>	60704,
		10649	=>	60705,
		10650	=>	60707,
		10651	=>	60709,
		10652	=>	60710,
		10653	=>	60712,
		10654	=>	60714,
		10655	=>	60715,
		10656	=>	60717,
		10657	=>	60719,
		10658	=>	60720,
		10659	=>	60722,
		10660	=>	60723,
		10661	=>	60725,
		10662	=>	60727,
		10663	=>	60728,
		10664	=>	60730,
		10665	=>	60732,
		10666	=>	60733,
		10667	=>	60735,
		10668	=>	60737,
		10669	=>	60738,
		10670	=>	60740,
		10671	=>	60741,
		10672	=>	60743,
		10673	=>	60745,
		10674	=>	60746,
		10675	=>	60748,
		10676	=>	60750,
		10677	=>	60751,
		10678	=>	60753,
		10679	=>	60755,
		10680	=>	60756,
		10681	=>	60758,
		10682	=>	60759,
		10683	=>	60761,
		10684	=>	60763,
		10685	=>	60764,
		10686	=>	60766,
		10687	=>	60768,
		10688	=>	60769,
		10689	=>	60771,
		10690	=>	60772,
		10691	=>	60774,
		10692	=>	60776,
		10693	=>	60777,
		10694	=>	60779,
		10695	=>	60781,
		10696	=>	60782,
		10697	=>	60784,
		10698	=>	60786,
		10699	=>	60787,
		10700	=>	60789,
		10701	=>	60790,
		10702	=>	60792,
		10703	=>	60794,
		10704	=>	60795,
		10705	=>	60797,
		10706	=>	60799,
		10707	=>	60800,
		10708	=>	60802,
		10709	=>	60803,
		10710	=>	60805,
		10711	=>	60807,
		10712	=>	60808,
		10713	=>	60810,
		10714	=>	60812,
		10715	=>	60813,
		10716	=>	60815,
		10717	=>	60816,
		10718	=>	60818,
		10719	=>	60820,
		10720	=>	60821,
		10721	=>	60823,
		10722	=>	60825,
		10723	=>	60826,
		10724	=>	60828,
		10725	=>	60829,
		10726	=>	60831,
		10727	=>	60833,
		10728	=>	60834,
		10729	=>	60836,
		10730	=>	60838,
		10731	=>	60839,
		10732	=>	60841,
		10733	=>	60842,
		10734	=>	60844,
		10735	=>	60846,
		10736	=>	60847,
		10737	=>	60849,
		10738	=>	60850,
		10739	=>	60852,
		10740	=>	60854,
		10741	=>	60855,
		10742	=>	60857,
		10743	=>	60859,
		10744	=>	60860,
		10745	=>	60862,
		10746	=>	60863,
		10747	=>	60865,
		10748	=>	60867,
		10749	=>	60868,
		10750	=>	60870,
		10751	=>	60872,
		10752	=>	60873,
		10753	=>	60875,
		10754	=>	60876,
		10755	=>	60878,
		10756	=>	60880,
		10757	=>	60881,
		10758	=>	60883,
		10759	=>	60884,
		10760	=>	60886,
		10761	=>	60888,
		10762	=>	60889,
		10763	=>	60891,
		10764	=>	60892,
		10765	=>	60894,
		10766	=>	60896,
		10767	=>	60897,
		10768	=>	60899,
		10769	=>	60901,
		10770	=>	60902,
		10771	=>	60904,
		10772	=>	60905,
		10773	=>	60907,
		10774	=>	60909,
		10775	=>	60910,
		10776	=>	60912,
		10777	=>	60913,
		10778	=>	60915,
		10779	=>	60917,
		10780	=>	60918,
		10781	=>	60920,
		10782	=>	60921,
		10783	=>	60923,
		10784	=>	60925,
		10785	=>	60926,
		10786	=>	60928,
		10787	=>	60929,
		10788	=>	60931,
		10789	=>	60933,
		10790	=>	60934,
		10791	=>	60936,
		10792	=>	60938,
		10793	=>	60939,
		10794	=>	60941,
		10795	=>	60942,
		10796	=>	60944,
		10797	=>	60946,
		10798	=>	60947,
		10799	=>	60949,
		10800	=>	60950,
		10801	=>	60952,
		10802	=>	60954,
		10803	=>	60955,
		10804	=>	60957,
		10805	=>	60958,
		10806	=>	60960,
		10807	=>	60962,
		10808	=>	60963,
		10809	=>	60965,
		10810	=>	60966,
		10811	=>	60968,
		10812	=>	60970,
		10813	=>	60971,
		10814	=>	60973,
		10815	=>	60974,
		10816	=>	60976,
		10817	=>	60978,
		10818	=>	60979,
		10819	=>	60981,
		10820	=>	60982,
		10821	=>	60984,
		10822	=>	60986,
		10823	=>	60987,
		10824	=>	60989,
		10825	=>	60990,
		10826	=>	60992,
		10827	=>	60994,
		10828	=>	60995,
		10829	=>	60997,
		10830	=>	60998,
		10831	=>	61000,
		10832	=>	61002,
		10833	=>	61003,
		10834	=>	61005,
		10835	=>	61006,
		10836	=>	61008,
		10837	=>	61009,
		10838	=>	61011,
		10839	=>	61013,
		10840	=>	61014,
		10841	=>	61016,
		10842	=>	61017,
		10843	=>	61019,
		10844	=>	61021,
		10845	=>	61022,
		10846	=>	61024,
		10847	=>	61025,
		10848	=>	61027,
		10849	=>	61029,
		10850	=>	61030,
		10851	=>	61032,
		10852	=>	61033,
		10853	=>	61035,
		10854	=>	61037,
		10855	=>	61038,
		10856	=>	61040,
		10857	=>	61041,
		10858	=>	61043,
		10859	=>	61044,
		10860	=>	61046,
		10861	=>	61048,
		10862	=>	61049,
		10863	=>	61051,
		10864	=>	61052,
		10865	=>	61054,
		10866	=>	61056,
		10867	=>	61057,
		10868	=>	61059,
		10869	=>	61060,
		10870	=>	61062,
		10871	=>	61063,
		10872	=>	61065,
		10873	=>	61067,
		10874	=>	61068,
		10875	=>	61070,
		10876	=>	61071,
		10877	=>	61073,
		10878	=>	61075,
		10879	=>	61076,
		10880	=>	61078,
		10881	=>	61079,
		10882	=>	61081,
		10883	=>	61082,
		10884	=>	61084,
		10885	=>	61086,
		10886	=>	61087,
		10887	=>	61089,
		10888	=>	61090,
		10889	=>	61092,
		10890	=>	61094,
		10891	=>	61095,
		10892	=>	61097,
		10893	=>	61098,
		10894	=>	61100,
		10895	=>	61101,
		10896	=>	61103,
		10897	=>	61105,
		10898	=>	61106,
		10899	=>	61108,
		10900	=>	61109,
		10901	=>	61111,
		10902	=>	61112,
		10903	=>	61114,
		10904	=>	61116,
		10905	=>	61117,
		10906	=>	61119,
		10907	=>	61120,
		10908	=>	61122,
		10909	=>	61123,
		10910	=>	61125,
		10911	=>	61127,
		10912	=>	61128,
		10913	=>	61130,
		10914	=>	61131,
		10915	=>	61133,
		10916	=>	61135,
		10917	=>	61136,
		10918	=>	61138,
		10919	=>	61139,
		10920	=>	61141,
		10921	=>	61142,
		10922	=>	61144,
		10923	=>	61146,
		10924	=>	61147,
		10925	=>	61149,
		10926	=>	61150,
		10927	=>	61152,
		10928	=>	61153,
		10929	=>	61155,
		10930	=>	61156,
		10931	=>	61158,
		10932	=>	61160,
		10933	=>	61161,
		10934	=>	61163,
		10935	=>	61164,
		10936	=>	61166,
		10937	=>	61167,
		10938	=>	61169,
		10939	=>	61171,
		10940	=>	61172,
		10941	=>	61174,
		10942	=>	61175,
		10943	=>	61177,
		10944	=>	61178,
		10945	=>	61180,
		10946	=>	61182,
		10947	=>	61183,
		10948	=>	61185,
		10949	=>	61186,
		10950	=>	61188,
		10951	=>	61189,
		10952	=>	61191,
		10953	=>	61193,
		10954	=>	61194,
		10955	=>	61196,
		10956	=>	61197,
		10957	=>	61199,
		10958	=>	61200,
		10959	=>	61202,
		10960	=>	61203,
		10961	=>	61205,
		10962	=>	61207,
		10963	=>	61208,
		10964	=>	61210,
		10965	=>	61211,
		10966	=>	61213,
		10967	=>	61214,
		10968	=>	61216,
		10969	=>	61217,
		10970	=>	61219,
		10971	=>	61221,
		10972	=>	61222,
		10973	=>	61224,
		10974	=>	61225,
		10975	=>	61227,
		10976	=>	61228,
		10977	=>	61230,
		10978	=>	61232,
		10979	=>	61233,
		10980	=>	61235,
		10981	=>	61236,
		10982	=>	61238,
		10983	=>	61239,
		10984	=>	61241,
		10985	=>	61242,
		10986	=>	61244,
		10987	=>	61246,
		10988	=>	61247,
		10989	=>	61249,
		10990	=>	61250,
		10991	=>	61252,
		10992	=>	61253,
		10993	=>	61255,
		10994	=>	61256,
		10995	=>	61258,
		10996	=>	61259,
		10997	=>	61261,
		10998	=>	61263,
		10999	=>	61264,
		11000	=>	61266,
		11001	=>	61267,
		11002	=>	61269,
		11003	=>	61270,
		11004	=>	61272,
		11005	=>	61273,
		11006	=>	61275,
		11007	=>	61277,
		11008	=>	61278,
		11009	=>	61280,
		11010	=>	61281,
		11011	=>	61283,
		11012	=>	61284,
		11013	=>	61286,
		11014	=>	61287,
		11015	=>	61289,
		11016	=>	61290,
		11017	=>	61292,
		11018	=>	61294,
		11019	=>	61295,
		11020	=>	61297,
		11021	=>	61298,
		11022	=>	61300,
		11023	=>	61301,
		11024	=>	61303,
		11025	=>	61304,
		11026	=>	61306,
		11027	=>	61307,
		11028	=>	61309,
		11029	=>	61311,
		11030	=>	61312,
		11031	=>	61314,
		11032	=>	61315,
		11033	=>	61317,
		11034	=>	61318,
		11035	=>	61320,
		11036	=>	61321,
		11037	=>	61323,
		11038	=>	61324,
		11039	=>	61326,
		11040	=>	61327,
		11041	=>	61329,
		11042	=>	61331,
		11043	=>	61332,
		11044	=>	61334,
		11045	=>	61335,
		11046	=>	61337,
		11047	=>	61338,
		11048	=>	61340,
		11049	=>	61341,
		11050	=>	61343,
		11051	=>	61344,
		11052	=>	61346,
		11053	=>	61347,
		11054	=>	61349,
		11055	=>	61351,
		11056	=>	61352,
		11057	=>	61354,
		11058	=>	61355,
		11059	=>	61357,
		11060	=>	61358,
		11061	=>	61360,
		11062	=>	61361,
		11063	=>	61363,
		11064	=>	61364,
		11065	=>	61366,
		11066	=>	61367,
		11067	=>	61369,
		11068	=>	61371,
		11069	=>	61372,
		11070	=>	61374,
		11071	=>	61375,
		11072	=>	61377,
		11073	=>	61378,
		11074	=>	61380,
		11075	=>	61381,
		11076	=>	61383,
		11077	=>	61384,
		11078	=>	61386,
		11079	=>	61387,
		11080	=>	61389,
		11081	=>	61390,
		11082	=>	61392,
		11083	=>	61393,
		11084	=>	61395,
		11085	=>	61397,
		11086	=>	61398,
		11087	=>	61400,
		11088	=>	61401,
		11089	=>	61403,
		11090	=>	61404,
		11091	=>	61406,
		11092	=>	61407,
		11093	=>	61409,
		11094	=>	61410,
		11095	=>	61412,
		11096	=>	61413,
		11097	=>	61415,
		11098	=>	61416,
		11099	=>	61418,
		11100	=>	61419,
		11101	=>	61421,
		11102	=>	61422,
		11103	=>	61424,
		11104	=>	61426,
		11105	=>	61427,
		11106	=>	61429,
		11107	=>	61430,
		11108	=>	61432,
		11109	=>	61433,
		11110	=>	61435,
		11111	=>	61436,
		11112	=>	61438,
		11113	=>	61439,
		11114	=>	61441,
		11115	=>	61442,
		11116	=>	61444,
		11117	=>	61445,
		11118	=>	61447,
		11119	=>	61448,
		11120	=>	61450,
		11121	=>	61451,
		11122	=>	61453,
		11123	=>	61454,
		11124	=>	61456,
		11125	=>	61457,
		11126	=>	61459,
		11127	=>	61460,
		11128	=>	61462,
		11129	=>	61464,
		11130	=>	61465,
		11131	=>	61467,
		11132	=>	61468,
		11133	=>	61470,
		11134	=>	61471,
		11135	=>	61473,
		11136	=>	61474,
		11137	=>	61476,
		11138	=>	61477,
		11139	=>	61479,
		11140	=>	61480,
		11141	=>	61482,
		11142	=>	61483,
		11143	=>	61485,
		11144	=>	61486,
		11145	=>	61488,
		11146	=>	61489,
		11147	=>	61491,
		11148	=>	61492,
		11149	=>	61494,
		11150	=>	61495,
		11151	=>	61497,
		11152	=>	61498,
		11153	=>	61500,
		11154	=>	61501,
		11155	=>	61503,
		11156	=>	61504,
		11157	=>	61506,
		11158	=>	61507,
		11159	=>	61509,
		11160	=>	61510,
		11161	=>	61512,
		11162	=>	61513,
		11163	=>	61515,
		11164	=>	61516,
		11165	=>	61518,
		11166	=>	61519,
		11167	=>	61521,
		11168	=>	61522,
		11169	=>	61524,
		11170	=>	61525,
		11171	=>	61527,
		11172	=>	61528,
		11173	=>	61530,
		11174	=>	61531,
		11175	=>	61533,
		11176	=>	61535,
		11177	=>	61536,
		11178	=>	61538,
		11179	=>	61539,
		11180	=>	61541,
		11181	=>	61542,
		11182	=>	61544,
		11183	=>	61545,
		11184	=>	61547,
		11185	=>	61548,
		11186	=>	61550,
		11187	=>	61551,
		11188	=>	61553,
		11189	=>	61554,
		11190	=>	61556,
		11191	=>	61557,
		11192	=>	61559,
		11193	=>	61560,
		11194	=>	61562,
		11195	=>	61563,
		11196	=>	61565,
		11197	=>	61566,
		11198	=>	61568,
		11199	=>	61569,
		11200	=>	61571,
		11201	=>	61572,
		11202	=>	61574,
		11203	=>	61575,
		11204	=>	61577,
		11205	=>	61578,
		11206	=>	61580,
		11207	=>	61581,
		11208	=>	61583,
		11209	=>	61584,
		11210	=>	61585,
		11211	=>	61587,
		11212	=>	61588,
		11213	=>	61590,
		11214	=>	61591,
		11215	=>	61593,
		11216	=>	61594,
		11217	=>	61596,
		11218	=>	61597,
		11219	=>	61599,
		11220	=>	61600,
		11221	=>	61602,
		11222	=>	61603,
		11223	=>	61605,
		11224	=>	61606,
		11225	=>	61608,
		11226	=>	61609,
		11227	=>	61611,
		11228	=>	61612,
		11229	=>	61614,
		11230	=>	61615,
		11231	=>	61617,
		11232	=>	61618,
		11233	=>	61620,
		11234	=>	61621,
		11235	=>	61623,
		11236	=>	61624,
		11237	=>	61626,
		11238	=>	61627,
		11239	=>	61629,
		11240	=>	61630,
		11241	=>	61632,
		11242	=>	61633,
		11243	=>	61635,
		11244	=>	61636,
		11245	=>	61638,
		11246	=>	61639,
		11247	=>	61641,
		11248	=>	61642,
		11249	=>	61644,
		11250	=>	61645,
		11251	=>	61647,
		11252	=>	61648,
		11253	=>	61650,
		11254	=>	61651,
		11255	=>	61653,
		11256	=>	61654,
		11257	=>	61655,
		11258	=>	61657,
		11259	=>	61658,
		11260	=>	61660,
		11261	=>	61661,
		11262	=>	61663,
		11263	=>	61664,
		11264	=>	61666,
		11265	=>	61667,
		11266	=>	61669,
		11267	=>	61670,
		11268	=>	61672,
		11269	=>	61673,
		11270	=>	61675,
		11271	=>	61676,
		11272	=>	61678,
		11273	=>	61679,
		11274	=>	61681,
		11275	=>	61682,
		11276	=>	61684,
		11277	=>	61685,
		11278	=>	61687,
		11279	=>	61688,
		11280	=>	61690,
		11281	=>	61691,
		11282	=>	61692,
		11283	=>	61694,
		11284	=>	61695,
		11285	=>	61697,
		11286	=>	61698,
		11287	=>	61700,
		11288	=>	61701,
		11289	=>	61703,
		11290	=>	61704,
		11291	=>	61706,
		11292	=>	61707,
		11293	=>	61709,
		11294	=>	61710,
		11295	=>	61712,
		11296	=>	61713,
		11297	=>	61715,
		11298	=>	61716,
		11299	=>	61718,
		11300	=>	61719,
		11301	=>	61720,
		11302	=>	61722,
		11303	=>	61723,
		11304	=>	61725,
		11305	=>	61726,
		11306	=>	61728,
		11307	=>	61729,
		11308	=>	61731,
		11309	=>	61732,
		11310	=>	61734,
		11311	=>	61735,
		11312	=>	61737,
		11313	=>	61738,
		11314	=>	61740,
		11315	=>	61741,
		11316	=>	61743,
		11317	=>	61744,
		11318	=>	61745,
		11319	=>	61747,
		11320	=>	61748,
		11321	=>	61750,
		11322	=>	61751,
		11323	=>	61753,
		11324	=>	61754,
		11325	=>	61756,
		11326	=>	61757,
		11327	=>	61759,
		11328	=>	61760,
		11329	=>	61762,
		11330	=>	61763,
		11331	=>	61764,
		11332	=>	61766,
		11333	=>	61767,
		11334	=>	61769,
		11335	=>	61770,
		11336	=>	61772,
		11337	=>	61773,
		11338	=>	61775,
		11339	=>	61776,
		11340	=>	61778,
		11341	=>	61779,
		11342	=>	61781,
		11343	=>	61782,
		11344	=>	61783,
		11345	=>	61785,
		11346	=>	61786,
		11347	=>	61788,
		11348	=>	61789,
		11349	=>	61791,
		11350	=>	61792,
		11351	=>	61794,
		11352	=>	61795,
		11353	=>	61797,
		11354	=>	61798,
		11355	=>	61800,
		11356	=>	61801,
		11357	=>	61802,
		11358	=>	61804,
		11359	=>	61805,
		11360	=>	61807,
		11361	=>	61808,
		11362	=>	61810,
		11363	=>	61811,
		11364	=>	61813,
		11365	=>	61814,
		11366	=>	61816,
		11367	=>	61817,
		11368	=>	61818,
		11369	=>	61820,
		11370	=>	61821,
		11371	=>	61823,
		11372	=>	61824,
		11373	=>	61826,
		11374	=>	61827,
		11375	=>	61829,
		11376	=>	61830,
		11377	=>	61831,
		11378	=>	61833,
		11379	=>	61834,
		11380	=>	61836,
		11381	=>	61837,
		11382	=>	61839,
		11383	=>	61840,
		11384	=>	61842,
		11385	=>	61843,
		11386	=>	61845,
		11387	=>	61846,
		11388	=>	61847,
		11389	=>	61849,
		11390	=>	61850,
		11391	=>	61852,
		11392	=>	61853,
		11393	=>	61855,
		11394	=>	61856,
		11395	=>	61858,
		11396	=>	61859,
		11397	=>	61860,
		11398	=>	61862,
		11399	=>	61863,
		11400	=>	61865,
		11401	=>	61866,
		11402	=>	61868,
		11403	=>	61869,
		11404	=>	61871,
		11405	=>	61872,
		11406	=>	61873,
		11407	=>	61875,
		11408	=>	61876,
		11409	=>	61878,
		11410	=>	61879,
		11411	=>	61881,
		11412	=>	61882,
		11413	=>	61884,
		11414	=>	61885,
		11415	=>	61886,
		11416	=>	61888,
		11417	=>	61889,
		11418	=>	61891,
		11419	=>	61892,
		11420	=>	61894,
		11421	=>	61895,
		11422	=>	61897,
		11423	=>	61898,
		11424	=>	61899,
		11425	=>	61901,
		11426	=>	61902,
		11427	=>	61904,
		11428	=>	61905,
		11429	=>	61907,
		11430	=>	61908,
		11431	=>	61909,
		11432	=>	61911,
		11433	=>	61912,
		11434	=>	61914,
		11435	=>	61915,
		11436	=>	61917,
		11437	=>	61918,
		11438	=>	61920,
		11439	=>	61921,
		11440	=>	61922,
		11441	=>	61924,
		11442	=>	61925,
		11443	=>	61927,
		11444	=>	61928,
		11445	=>	61930,
		11446	=>	61931,
		11447	=>	61932,
		11448	=>	61934,
		11449	=>	61935,
		11450	=>	61937,
		11451	=>	61938,
		11452	=>	61940,
		11453	=>	61941,
		11454	=>	61942,
		11455	=>	61944,
		11456	=>	61945,
		11457	=>	61947,
		11458	=>	61948,
		11459	=>	61950,
		11460	=>	61951,
		11461	=>	61952,
		11462	=>	61954,
		11463	=>	61955,
		11464	=>	61957,
		11465	=>	61958,
		11466	=>	61960,
		11467	=>	61961,
		11468	=>	61962,
		11469	=>	61964,
		11470	=>	61965,
		11471	=>	61967,
		11472	=>	61968,
		11473	=>	61970,
		11474	=>	61971,
		11475	=>	61972,
		11476	=>	61974,
		11477	=>	61975,
		11478	=>	61977,
		11479	=>	61978,
		11480	=>	61980,
		11481	=>	61981,
		11482	=>	61982,
		11483	=>	61984,
		11484	=>	61985,
		11485	=>	61987,
		11486	=>	61988,
		11487	=>	61989,
		11488	=>	61991,
		11489	=>	61992,
		11490	=>	61994,
		11491	=>	61995,
		11492	=>	61997,
		11493	=>	61998,
		11494	=>	61999,
		11495	=>	62001,
		11496	=>	62002,
		11497	=>	62004,
		11498	=>	62005,
		11499	=>	62007,
		11500	=>	62008,
		11501	=>	62009,
		11502	=>	62011,
		11503	=>	62012,
		11504	=>	62014,
		11505	=>	62015,
		11506	=>	62016,
		11507	=>	62018,
		11508	=>	62019,
		11509	=>	62021,
		11510	=>	62022,
		11511	=>	62024,
		11512	=>	62025,
		11513	=>	62026,
		11514	=>	62028,
		11515	=>	62029,
		11516	=>	62031,
		11517	=>	62032,
		11518	=>	62033,
		11519	=>	62035,
		11520	=>	62036,
		11521	=>	62038,
		11522	=>	62039,
		11523	=>	62040,
		11524	=>	62042,
		11525	=>	62043,
		11526	=>	62045,
		11527	=>	62046,
		11528	=>	62048,
		11529	=>	62049,
		11530	=>	62050,
		11531	=>	62052,
		11532	=>	62053,
		11533	=>	62055,
		11534	=>	62056,
		11535	=>	62057,
		11536	=>	62059,
		11537	=>	62060,
		11538	=>	62062,
		11539	=>	62063,
		11540	=>	62064,
		11541	=>	62066,
		11542	=>	62067,
		11543	=>	62069,
		11544	=>	62070,
		11545	=>	62071,
		11546	=>	62073,
		11547	=>	62074,
		11548	=>	62076,
		11549	=>	62077,
		11550	=>	62078,
		11551	=>	62080,
		11552	=>	62081,
		11553	=>	62083,
		11554	=>	62084,
		11555	=>	62085,
		11556	=>	62087,
		11557	=>	62088,
		11558	=>	62090,
		11559	=>	62091,
		11560	=>	62093,
		11561	=>	62094,
		11562	=>	62095,
		11563	=>	62097,
		11564	=>	62098,
		11565	=>	62100,
		11566	=>	62101,
		11567	=>	62102,
		11568	=>	62104,
		11569	=>	62105,
		11570	=>	62107,
		11571	=>	62108,
		11572	=>	62109,
		11573	=>	62111,
		11574	=>	62112,
		11575	=>	62114,
		11576	=>	62115,
		11577	=>	62116,
		11578	=>	62118,
		11579	=>	62119,
		11580	=>	62120,
		11581	=>	62122,
		11582	=>	62123,
		11583	=>	62125,
		11584	=>	62126,
		11585	=>	62127,
		11586	=>	62129,
		11587	=>	62130,
		11588	=>	62132,
		11589	=>	62133,
		11590	=>	62134,
		11591	=>	62136,
		11592	=>	62137,
		11593	=>	62139,
		11594	=>	62140,
		11595	=>	62141,
		11596	=>	62143,
		11597	=>	62144,
		11598	=>	62146,
		11599	=>	62147,
		11600	=>	62148,
		11601	=>	62150,
		11602	=>	62151,
		11603	=>	62153,
		11604	=>	62154,
		11605	=>	62155,
		11606	=>	62157,
		11607	=>	62158,
		11608	=>	62159,
		11609	=>	62161,
		11610	=>	62162,
		11611	=>	62164,
		11612	=>	62165,
		11613	=>	62166,
		11614	=>	62168,
		11615	=>	62169,
		11616	=>	62171,
		11617	=>	62172,
		11618	=>	62173,
		11619	=>	62175,
		11620	=>	62176,
		11621	=>	62178,
		11622	=>	62179,
		11623	=>	62180,
		11624	=>	62182,
		11625	=>	62183,
		11626	=>	62184,
		11627	=>	62186,
		11628	=>	62187,
		11629	=>	62189,
		11630	=>	62190,
		11631	=>	62191,
		11632	=>	62193,
		11633	=>	62194,
		11634	=>	62195,
		11635	=>	62197,
		11636	=>	62198,
		11637	=>	62200,
		11638	=>	62201,
		11639	=>	62202,
		11640	=>	62204,
		11641	=>	62205,
		11642	=>	62207,
		11643	=>	62208,
		11644	=>	62209,
		11645	=>	62211,
		11646	=>	62212,
		11647	=>	62213,
		11648	=>	62215,
		11649	=>	62216,
		11650	=>	62218,
		11651	=>	62219,
		11652	=>	62220,
		11653	=>	62222,
		11654	=>	62223,
		11655	=>	62224,
		11656	=>	62226,
		11657	=>	62227,
		11658	=>	62229,
		11659	=>	62230,
		11660	=>	62231,
		11661	=>	62233,
		11662	=>	62234,
		11663	=>	62235,
		11664	=>	62237,
		11665	=>	62238,
		11666	=>	62240,
		11667	=>	62241,
		11668	=>	62242,
		11669	=>	62244,
		11670	=>	62245,
		11671	=>	62246,
		11672	=>	62248,
		11673	=>	62249,
		11674	=>	62251,
		11675	=>	62252,
		11676	=>	62253,
		11677	=>	62255,
		11678	=>	62256,
		11679	=>	62257,
		11680	=>	62259,
		11681	=>	62260,
		11682	=>	62262,
		11683	=>	62263,
		11684	=>	62264,
		11685	=>	62266,
		11686	=>	62267,
		11687	=>	62268,
		11688	=>	62270,
		11689	=>	62271,
		11690	=>	62272,
		11691	=>	62274,
		11692	=>	62275,
		11693	=>	62277,
		11694	=>	62278,
		11695	=>	62279,
		11696	=>	62281,
		11697	=>	62282,
		11698	=>	62283,
		11699	=>	62285,
		11700	=>	62286,
		11701	=>	62287,
		11702	=>	62289,
		11703	=>	62290,
		11704	=>	62292,
		11705	=>	62293,
		11706	=>	62294,
		11707	=>	62296,
		11708	=>	62297,
		11709	=>	62298,
		11710	=>	62300,
		11711	=>	62301,
		11712	=>	62302,
		11713	=>	62304,
		11714	=>	62305,
		11715	=>	62307,
		11716	=>	62308,
		11717	=>	62309,
		11718	=>	62311,
		11719	=>	62312,
		11720	=>	62313,
		11721	=>	62315,
		11722	=>	62316,
		11723	=>	62317,
		11724	=>	62319,
		11725	=>	62320,
		11726	=>	62321,
		11727	=>	62323,
		11728	=>	62324,
		11729	=>	62326,
		11730	=>	62327,
		11731	=>	62328,
		11732	=>	62330,
		11733	=>	62331,
		11734	=>	62332,
		11735	=>	62334,
		11736	=>	62335,
		11737	=>	62336,
		11738	=>	62338,
		11739	=>	62339,
		11740	=>	62340,
		11741	=>	62342,
		11742	=>	62343,
		11743	=>	62344,
		11744	=>	62346,
		11745	=>	62347,
		11746	=>	62349,
		11747	=>	62350,
		11748	=>	62351,
		11749	=>	62353,
		11750	=>	62354,
		11751	=>	62355,
		11752	=>	62357,
		11753	=>	62358,
		11754	=>	62359,
		11755	=>	62361,
		11756	=>	62362,
		11757	=>	62363,
		11758	=>	62365,
		11759	=>	62366,
		11760	=>	62367,
		11761	=>	62369,
		11762	=>	62370,
		11763	=>	62371,
		11764	=>	62373,
		11765	=>	62374,
		11766	=>	62376,
		11767	=>	62377,
		11768	=>	62378,
		11769	=>	62380,
		11770	=>	62381,
		11771	=>	62382,
		11772	=>	62384,
		11773	=>	62385,
		11774	=>	62386,
		11775	=>	62388,
		11776	=>	62389,
		11777	=>	62390,
		11778	=>	62392,
		11779	=>	62393,
		11780	=>	62394,
		11781	=>	62396,
		11782	=>	62397,
		11783	=>	62398,
		11784	=>	62400,
		11785	=>	62401,
		11786	=>	62402,
		11787	=>	62404,
		11788	=>	62405,
		11789	=>	62406,
		11790	=>	62408,
		11791	=>	62409,
		11792	=>	62410,
		11793	=>	62412,
		11794	=>	62413,
		11795	=>	62414,
		11796	=>	62416,
		11797	=>	62417,
		11798	=>	62418,
		11799	=>	62420,
		11800	=>	62421,
		11801	=>	62422,
		11802	=>	62424,
		11803	=>	62425,
		11804	=>	62426,
		11805	=>	62428,
		11806	=>	62429,
		11807	=>	62430,
		11808	=>	62432,
		11809	=>	62433,
		11810	=>	62434,
		11811	=>	62436,
		11812	=>	62437,
		11813	=>	62438,
		11814	=>	62440,
		11815	=>	62441,
		11816	=>	62442,
		11817	=>	62444,
		11818	=>	62445,
		11819	=>	62446,
		11820	=>	62448,
		11821	=>	62449,
		11822	=>	62450,
		11823	=>	62452,
		11824	=>	62453,
		11825	=>	62454,
		11826	=>	62456,
		11827	=>	62457,
		11828	=>	62458,
		11829	=>	62460,
		11830	=>	62461,
		11831	=>	62462,
		11832	=>	62464,
		11833	=>	62465,
		11834	=>	62466,
		11835	=>	62468,
		11836	=>	62469,
		11837	=>	62470,
		11838	=>	62472,
		11839	=>	62473,
		11840	=>	62474,
		11841	=>	62476,
		11842	=>	62477,
		11843	=>	62478,
		11844	=>	62480,
		11845	=>	62481,
		11846	=>	62482,
		11847	=>	62484,
		11848	=>	62485,
		11849	=>	62486,
		11850	=>	62488,
		11851	=>	62489,
		11852	=>	62490,
		11853	=>	62492,
		11854	=>	62493,
		11855	=>	62494,
		11856	=>	62496,
		11857	=>	62497,
		11858	=>	62498,
		11859	=>	62500,
		11860	=>	62501,
		11861	=>	62502,
		11862	=>	62503,
		11863	=>	62505,
		11864	=>	62506,
		11865	=>	62507,
		11866	=>	62509,
		11867	=>	62510,
		11868	=>	62511,
		11869	=>	62513,
		11870	=>	62514,
		11871	=>	62515,
		11872	=>	62517,
		11873	=>	62518,
		11874	=>	62519,
		11875	=>	62521,
		11876	=>	62522,
		11877	=>	62523,
		11878	=>	62525,
		11879	=>	62526,
		11880	=>	62527,
		11881	=>	62529,
		11882	=>	62530,
		11883	=>	62531,
		11884	=>	62532,
		11885	=>	62534,
		11886	=>	62535,
		11887	=>	62536,
		11888	=>	62538,
		11889	=>	62539,
		11890	=>	62540,
		11891	=>	62542,
		11892	=>	62543,
		11893	=>	62544,
		11894	=>	62546,
		11895	=>	62547,
		11896	=>	62548,
		11897	=>	62549,
		11898	=>	62551,
		11899	=>	62552,
		11900	=>	62553,
		11901	=>	62555,
		11902	=>	62556,
		11903	=>	62557,
		11904	=>	62559,
		11905	=>	62560,
		11906	=>	62561,
		11907	=>	62563,
		11908	=>	62564,
		11909	=>	62565,
		11910	=>	62567,
		11911	=>	62568,
		11912	=>	62569,
		11913	=>	62570,
		11914	=>	62572,
		11915	=>	62573,
		11916	=>	62574,
		11917	=>	62576,
		11918	=>	62577,
		11919	=>	62578,
		11920	=>	62580,
		11921	=>	62581,
		11922	=>	62582,
		11923	=>	62583,
		11924	=>	62585,
		11925	=>	62586,
		11926	=>	62587,
		11927	=>	62589,
		11928	=>	62590,
		11929	=>	62591,
		11930	=>	62593,
		11931	=>	62594,
		11932	=>	62595,
		11933	=>	62596,
		11934	=>	62598,
		11935	=>	62599,
		11936	=>	62600,
		11937	=>	62602,
		11938	=>	62603,
		11939	=>	62604,
		11940	=>	62606,
		11941	=>	62607,
		11942	=>	62608,
		11943	=>	62609,
		11944	=>	62611,
		11945	=>	62612,
		11946	=>	62613,
		11947	=>	62615,
		11948	=>	62616,
		11949	=>	62617,
		11950	=>	62619,
		11951	=>	62620,
		11952	=>	62621,
		11953	=>	62622,
		11954	=>	62624,
		11955	=>	62625,
		11956	=>	62626,
		11957	=>	62628,
		11958	=>	62629,
		11959	=>	62630,
		11960	=>	62631,
		11961	=>	62633,
		11962	=>	62634,
		11963	=>	62635,
		11964	=>	62637,
		11965	=>	62638,
		11966	=>	62639,
		11967	=>	62641,
		11968	=>	62642,
		11969	=>	62643,
		11970	=>	62644,
		11971	=>	62646,
		11972	=>	62647,
		11973	=>	62648,
		11974	=>	62650,
		11975	=>	62651,
		11976	=>	62652,
		11977	=>	62653,
		11978	=>	62655,
		11979	=>	62656,
		11980	=>	62657,
		11981	=>	62659,
		11982	=>	62660,
		11983	=>	62661,
		11984	=>	62662,
		11985	=>	62664,
		11986	=>	62665,
		11987	=>	62666,
		11988	=>	62668,
		11989	=>	62669,
		11990	=>	62670,
		11991	=>	62671,
		11992	=>	62673,
		11993	=>	62674,
		11994	=>	62675,
		11995	=>	62677,
		11996	=>	62678,
		11997	=>	62679,
		11998	=>	62680,
		11999	=>	62682,
		12000	=>	62683,
		12001	=>	62684,
		12002	=>	62686,
		12003	=>	62687,
		12004	=>	62688,
		12005	=>	62689,
		12006	=>	62691,
		12007	=>	62692,
		12008	=>	62693,
		12009	=>	62695,
		12010	=>	62696,
		12011	=>	62697,
		12012	=>	62698,
		12013	=>	62700,
		12014	=>	62701,
		12015	=>	62702,
		12016	=>	62703,
		12017	=>	62705,
		12018	=>	62706,
		12019	=>	62707,
		12020	=>	62709,
		12021	=>	62710,
		12022	=>	62711,
		12023	=>	62712,
		12024	=>	62714,
		12025	=>	62715,
		12026	=>	62716,
		12027	=>	62717,
		12028	=>	62719,
		12029	=>	62720,
		12030	=>	62721,
		12031	=>	62723,
		12032	=>	62724,
		12033	=>	62725,
		12034	=>	62726,
		12035	=>	62728,
		12036	=>	62729,
		12037	=>	62730,
		12038	=>	62732,
		12039	=>	62733,
		12040	=>	62734,
		12041	=>	62735,
		12042	=>	62737,
		12043	=>	62738,
		12044	=>	62739,
		12045	=>	62740,
		12046	=>	62742,
		12047	=>	62743,
		12048	=>	62744,
		12049	=>	62745,
		12050	=>	62747,
		12051	=>	62748,
		12052	=>	62749,
		12053	=>	62751,
		12054	=>	62752,
		12055	=>	62753,
		12056	=>	62754,
		12057	=>	62756,
		12058	=>	62757,
		12059	=>	62758,
		12060	=>	62759,
		12061	=>	62761,
		12062	=>	62762,
		12063	=>	62763,
		12064	=>	62764,
		12065	=>	62766,
		12066	=>	62767,
		12067	=>	62768,
		12068	=>	62770,
		12069	=>	62771,
		12070	=>	62772,
		12071	=>	62773,
		12072	=>	62775,
		12073	=>	62776,
		12074	=>	62777,
		12075	=>	62778,
		12076	=>	62780,
		12077	=>	62781,
		12078	=>	62782,
		12079	=>	62783,
		12080	=>	62785,
		12081	=>	62786,
		12082	=>	62787,
		12083	=>	62788,
		12084	=>	62790,
		12085	=>	62791,
		12086	=>	62792,
		12087	=>	62793,
		12088	=>	62795,
		12089	=>	62796,
		12090	=>	62797,
		12091	=>	62799,
		12092	=>	62800,
		12093	=>	62801,
		12094	=>	62802,
		12095	=>	62804,
		12096	=>	62805,
		12097	=>	62806,
		12098	=>	62807,
		12099	=>	62809,
		12100	=>	62810,
		12101	=>	62811,
		12102	=>	62812,
		12103	=>	62814,
		12104	=>	62815,
		12105	=>	62816,
		12106	=>	62817,
		12107	=>	62819,
		12108	=>	62820,
		12109	=>	62821,
		12110	=>	62822,
		12111	=>	62824,
		12112	=>	62825,
		12113	=>	62826,
		12114	=>	62827,
		12115	=>	62829,
		12116	=>	62830,
		12117	=>	62831,
		12118	=>	62832,
		12119	=>	62834,
		12120	=>	62835,
		12121	=>	62836,
		12122	=>	62837,
		12123	=>	62839,
		12124	=>	62840,
		12125	=>	62841,
		12126	=>	62842,
		12127	=>	62844,
		12128	=>	62845,
		12129	=>	62846,
		12130	=>	62847,
		12131	=>	62849,
		12132	=>	62850,
		12133	=>	62851,
		12134	=>	62852,
		12135	=>	62854,
		12136	=>	62855,
		12137	=>	62856,
		12138	=>	62857,
		12139	=>	62859,
		12140	=>	62860,
		12141	=>	62861,
		12142	=>	62862,
		12143	=>	62863,
		12144	=>	62865,
		12145	=>	62866,
		12146	=>	62867,
		12147	=>	62868,
		12148	=>	62870,
		12149	=>	62871,
		12150	=>	62872,
		12151	=>	62873,
		12152	=>	62875,
		12153	=>	62876,
		12154	=>	62877,
		12155	=>	62878,
		12156	=>	62880,
		12157	=>	62881,
		12158	=>	62882,
		12159	=>	62883,
		12160	=>	62885,
		12161	=>	62886,
		12162	=>	62887,
		12163	=>	62888,
		12164	=>	62890,
		12165	=>	62891,
		12166	=>	62892,
		12167	=>	62893,
		12168	=>	62894,
		12169	=>	62896,
		12170	=>	62897,
		12171	=>	62898,
		12172	=>	62899,
		12173	=>	62901,
		12174	=>	62902,
		12175	=>	62903,
		12176	=>	62904,
		12177	=>	62906,
		12178	=>	62907,
		12179	=>	62908,
		12180	=>	62909,
		12181	=>	62910,
		12182	=>	62912,
		12183	=>	62913,
		12184	=>	62914,
		12185	=>	62915,
		12186	=>	62917,
		12187	=>	62918,
		12188	=>	62919,
		12189	=>	62920,
		12190	=>	62922,
		12191	=>	62923,
		12192	=>	62924,
		12193	=>	62925,
		12194	=>	62926,
		12195	=>	62928,
		12196	=>	62929,
		12197	=>	62930,
		12198	=>	62931,
		12199	=>	62933,
		12200	=>	62934,
		12201	=>	62935,
		12202	=>	62936,
		12203	=>	62938,
		12204	=>	62939,
		12205	=>	62940,
		12206	=>	62941,
		12207	=>	62942,
		12208	=>	62944,
		12209	=>	62945,
		12210	=>	62946,
		12211	=>	62947,
		12212	=>	62949,
		12213	=>	62950,
		12214	=>	62951,
		12215	=>	62952,
		12216	=>	62953,
		12217	=>	62955,
		12218	=>	62956,
		12219	=>	62957,
		12220	=>	62958,
		12221	=>	62960,
		12222	=>	62961,
		12223	=>	62962,
		12224	=>	62963,
		12225	=>	62964,
		12226	=>	62966,
		12227	=>	62967,
		12228	=>	62968,
		12229	=>	62969,
		12230	=>	62971,
		12231	=>	62972,
		12232	=>	62973,
		12233	=>	62974,
		12234	=>	62975,
		12235	=>	62977,
		12236	=>	62978,
		12237	=>	62979,
		12238	=>	62980,
		12239	=>	62981,
		12240	=>	62983,
		12241	=>	62984,
		12242	=>	62985,
		12243	=>	62986,
		12244	=>	62988,
		12245	=>	62989,
		12246	=>	62990,
		12247	=>	62991,
		12248	=>	62992,
		12249	=>	62994,
		12250	=>	62995,
		12251	=>	62996,
		12252	=>	62997,
		12253	=>	62998,
		12254	=>	63000,
		12255	=>	63001,
		12256	=>	63002,
		12257	=>	63003,
		12258	=>	63005,
		12259	=>	63006,
		12260	=>	63007,
		12261	=>	63008,
		12262	=>	63009,
		12263	=>	63011,
		12264	=>	63012,
		12265	=>	63013,
		12266	=>	63014,
		12267	=>	63015,
		12268	=>	63017,
		12269	=>	63018,
		12270	=>	63019,
		12271	=>	63020,
		12272	=>	63021,
		12273	=>	63023,
		12274	=>	63024,
		12275	=>	63025,
		12276	=>	63026,
		12277	=>	63027,
		12278	=>	63029,
		12279	=>	63030,
		12280	=>	63031,
		12281	=>	63032,
		12282	=>	63034,
		12283	=>	63035,
		12284	=>	63036,
		12285	=>	63037,
		12286	=>	63038,
		12287	=>	63040,
		12288	=>	63041,
		12289	=>	63042,
		12290	=>	63043,
		12291	=>	63044,
		12292	=>	63046,
		12293	=>	63047,
		12294	=>	63048,
		12295	=>	63049,
		12296	=>	63050,
		12297	=>	63052,
		12298	=>	63053,
		12299	=>	63054,
		12300	=>	63055,
		12301	=>	63056,
		12302	=>	63058,
		12303	=>	63059,
		12304	=>	63060,
		12305	=>	63061,
		12306	=>	63062,
		12307	=>	63064,
		12308	=>	63065,
		12309	=>	63066,
		12310	=>	63067,
		12311	=>	63068,
		12312	=>	63069,
		12313	=>	63071,
		12314	=>	63072,
		12315	=>	63073,
		12316	=>	63074,
		12317	=>	63075,
		12318	=>	63077,
		12319	=>	63078,
		12320	=>	63079,
		12321	=>	63080,
		12322	=>	63081,
		12323	=>	63083,
		12324	=>	63084,
		12325	=>	63085,
		12326	=>	63086,
		12327	=>	63087,
		12328	=>	63089,
		12329	=>	63090,
		12330	=>	63091,
		12331	=>	63092,
		12332	=>	63093,
		12333	=>	63095,
		12334	=>	63096,
		12335	=>	63097,
		12336	=>	63098,
		12337	=>	63099,
		12338	=>	63100,
		12339	=>	63102,
		12340	=>	63103,
		12341	=>	63104,
		12342	=>	63105,
		12343	=>	63106,
		12344	=>	63108,
		12345	=>	63109,
		12346	=>	63110,
		12347	=>	63111,
		12348	=>	63112,
		12349	=>	63114,
		12350	=>	63115,
		12351	=>	63116,
		12352	=>	63117,
		12353	=>	63118,
		12354	=>	63119,
		12355	=>	63121,
		12356	=>	63122,
		12357	=>	63123,
		12358	=>	63124,
		12359	=>	63125,
		12360	=>	63127,
		12361	=>	63128,
		12362	=>	63129,
		12363	=>	63130,
		12364	=>	63131,
		12365	=>	63132,
		12366	=>	63134,
		12367	=>	63135,
		12368	=>	63136,
		12369	=>	63137,
		12370	=>	63138,
		12371	=>	63140,
		12372	=>	63141,
		12373	=>	63142,
		12374	=>	63143,
		12375	=>	63144,
		12376	=>	63145,
		12377	=>	63147,
		12378	=>	63148,
		12379	=>	63149,
		12380	=>	63150,
		12381	=>	63151,
		12382	=>	63153,
		12383	=>	63154,
		12384	=>	63155,
		12385	=>	63156,
		12386	=>	63157,
		12387	=>	63158,
		12388	=>	63160,
		12389	=>	63161,
		12390	=>	63162,
		12391	=>	63163,
		12392	=>	63164,
		12393	=>	63165,
		12394	=>	63167,
		12395	=>	63168,
		12396	=>	63169,
		12397	=>	63170,
		12398	=>	63171,
		12399	=>	63172,
		12400	=>	63174,
		12401	=>	63175,
		12402	=>	63176,
		12403	=>	63177,
		12404	=>	63178,
		12405	=>	63179,
		12406	=>	63181,
		12407	=>	63182,
		12408	=>	63183,
		12409	=>	63184,
		12410	=>	63185,
		12411	=>	63186,
		12412	=>	63188,
		12413	=>	63189,
		12414	=>	63190,
		12415	=>	63191,
		12416	=>	63192,
		12417	=>	63193,
		12418	=>	63195,
		12419	=>	63196,
		12420	=>	63197,
		12421	=>	63198,
		12422	=>	63199,
		12423	=>	63200,
		12424	=>	63202,
		12425	=>	63203,
		12426	=>	63204,
		12427	=>	63205,
		12428	=>	63206,
		12429	=>	63207,
		12430	=>	63209,
		12431	=>	63210,
		12432	=>	63211,
		12433	=>	63212,
		12434	=>	63213,
		12435	=>	63214,
		12436	=>	63216,
		12437	=>	63217,
		12438	=>	63218,
		12439	=>	63219,
		12440	=>	63220,
		12441	=>	63221,
		12442	=>	63223,
		12443	=>	63224,
		12444	=>	63225,
		12445	=>	63226,
		12446	=>	63227,
		12447	=>	63228,
		12448	=>	63230,
		12449	=>	63231,
		12450	=>	63232,
		12451	=>	63233,
		12452	=>	63234,
		12453	=>	63235,
		12454	=>	63236,
		12455	=>	63238,
		12456	=>	63239,
		12457	=>	63240,
		12458	=>	63241,
		12459	=>	63242,
		12460	=>	63243,
		12461	=>	63245,
		12462	=>	63246,
		12463	=>	63247,
		12464	=>	63248,
		12465	=>	63249,
		12466	=>	63250,
		12467	=>	63251,
		12468	=>	63253,
		12469	=>	63254,
		12470	=>	63255,
		12471	=>	63256,
		12472	=>	63257,
		12473	=>	63258,
		12474	=>	63260,
		12475	=>	63261,
		12476	=>	63262,
		12477	=>	63263,
		12478	=>	63264,
		12479	=>	63265,
		12480	=>	63266,
		12481	=>	63268,
		12482	=>	63269,
		12483	=>	63270,
		12484	=>	63271,
		12485	=>	63272,
		12486	=>	63273,
		12487	=>	63274,
		12488	=>	63276,
		12489	=>	63277,
		12490	=>	63278,
		12491	=>	63279,
		12492	=>	63280,
		12493	=>	63281,
		12494	=>	63282,
		12495	=>	63284,
		12496	=>	63285,
		12497	=>	63286,
		12498	=>	63287,
		12499	=>	63288,
		12500	=>	63289,
		12501	=>	63290,
		12502	=>	63292,
		12503	=>	63293,
		12504	=>	63294,
		12505	=>	63295,
		12506	=>	63296,
		12507	=>	63297,
		12508	=>	63298,
		12509	=>	63300,
		12510	=>	63301,
		12511	=>	63302,
		12512	=>	63303,
		12513	=>	63304,
		12514	=>	63305,
		12515	=>	63306,
		12516	=>	63308,
		12517	=>	63309,
		12518	=>	63310,
		12519	=>	63311,
		12520	=>	63312,
		12521	=>	63313,
		12522	=>	63314,
		12523	=>	63316,
		12524	=>	63317,
		12525	=>	63318,
		12526	=>	63319,
		12527	=>	63320,
		12528	=>	63321,
		12529	=>	63322,
		12530	=>	63323,
		12531	=>	63325,
		12532	=>	63326,
		12533	=>	63327,
		12534	=>	63328,
		12535	=>	63329,
		12536	=>	63330,
		12537	=>	63331,
		12538	=>	63333,
		12539	=>	63334,
		12540	=>	63335,
		12541	=>	63336,
		12542	=>	63337,
		12543	=>	63338,
		12544	=>	63339,
		12545	=>	63340,
		12546	=>	63342,
		12547	=>	63343,
		12548	=>	63344,
		12549	=>	63345,
		12550	=>	63346,
		12551	=>	63347,
		12552	=>	63348,
		12553	=>	63350,
		12554	=>	63351,
		12555	=>	63352,
		12556	=>	63353,
		12557	=>	63354,
		12558	=>	63355,
		12559	=>	63356,
		12560	=>	63357,
		12561	=>	63359,
		12562	=>	63360,
		12563	=>	63361,
		12564	=>	63362,
		12565	=>	63363,
		12566	=>	63364,
		12567	=>	63365,
		12568	=>	63366,
		12569	=>	63368,
		12570	=>	63369,
		12571	=>	63370,
		12572	=>	63371,
		12573	=>	63372,
		12574	=>	63373,
		12575	=>	63374,
		12576	=>	63375,
		12577	=>	63376,
		12578	=>	63378,
		12579	=>	63379,
		12580	=>	63380,
		12581	=>	63381,
		12582	=>	63382,
		12583	=>	63383,
		12584	=>	63384,
		12585	=>	63385,
		12586	=>	63387,
		12587	=>	63388,
		12588	=>	63389,
		12589	=>	63390,
		12590	=>	63391,
		12591	=>	63392,
		12592	=>	63393,
		12593	=>	63394,
		12594	=>	63396,
		12595	=>	63397,
		12596	=>	63398,
		12597	=>	63399,
		12598	=>	63400,
		12599	=>	63401,
		12600	=>	63402,
		12601	=>	63403,
		12602	=>	63404,
		12603	=>	63406,
		12604	=>	63407,
		12605	=>	63408,
		12606	=>	63409,
		12607	=>	63410,
		12608	=>	63411,
		12609	=>	63412,
		12610	=>	63413,
		12611	=>	63414,
		12612	=>	63416,
		12613	=>	63417,
		12614	=>	63418,
		12615	=>	63419,
		12616	=>	63420,
		12617	=>	63421,
		12618	=>	63422,
		12619	=>	63423,
		12620	=>	63424,
		12621	=>	63426,
		12622	=>	63427,
		12623	=>	63428,
		12624	=>	63429,
		12625	=>	63430,
		12626	=>	63431,
		12627	=>	63432,
		12628	=>	63433,
		12629	=>	63434,
		12630	=>	63436,
		12631	=>	63437,
		12632	=>	63438,
		12633	=>	63439,
		12634	=>	63440,
		12635	=>	63441,
		12636	=>	63442,
		12637	=>	63443,
		12638	=>	63444,
		12639	=>	63445,
		12640	=>	63447,
		12641	=>	63448,
		12642	=>	63449,
		12643	=>	63450,
		12644	=>	63451,
		12645	=>	63452,
		12646	=>	63453,
		12647	=>	63454,
		12648	=>	63455,
		12649	=>	63457,
		12650	=>	63458,
		12651	=>	63459,
		12652	=>	63460,
		12653	=>	63461,
		12654	=>	63462,
		12655	=>	63463,
		12656	=>	63464,
		12657	=>	63465,
		12658	=>	63466,
		12659	=>	63468,
		12660	=>	63469,
		12661	=>	63470,
		12662	=>	63471,
		12663	=>	63472,
		12664	=>	63473,
		12665	=>	63474,
		12666	=>	63475,
		12667	=>	63476,
		12668	=>	63477,
		12669	=>	63478,
		12670	=>	63480,
		12671	=>	63481,
		12672	=>	63482,
		12673	=>	63483,
		12674	=>	63484,
		12675	=>	63485,
		12676	=>	63486,
		12677	=>	63487,
		12678	=>	63488,
		12679	=>	63489,
		12680	=>	63491,
		12681	=>	63492,
		12682	=>	63493,
		12683	=>	63494,
		12684	=>	63495,
		12685	=>	63496,
		12686	=>	63497,
		12687	=>	63498,
		12688	=>	63499,
		12689	=>	63500,
		12690	=>	63501,
		12691	=>	63503,
		12692	=>	63504,
		12693	=>	63505,
		12694	=>	63506,
		12695	=>	63507,
		12696	=>	63508,
		12697	=>	63509,
		12698	=>	63510,
		12699	=>	63511,
		12700	=>	63512,
		12701	=>	63513,
		12702	=>	63514,
		12703	=>	63516,
		12704	=>	63517,
		12705	=>	63518,
		12706	=>	63519,
		12707	=>	63520,
		12708	=>	63521,
		12709	=>	63522,
		12710	=>	63523,
		12711	=>	63524,
		12712	=>	63525,
		12713	=>	63526,
		12714	=>	63527,
		12715	=>	63529,
		12716	=>	63530,
		12717	=>	63531,
		12718	=>	63532,
		12719	=>	63533,
		12720	=>	63534,
		12721	=>	63535,
		12722	=>	63536,
		12723	=>	63537,
		12724	=>	63538,
		12725	=>	63539,
		12726	=>	63540,
		12727	=>	63542,
		12728	=>	63543,
		12729	=>	63544,
		12730	=>	63545,
		12731	=>	63546,
		12732	=>	63547,
		12733	=>	63548,
		12734	=>	63549,
		12735	=>	63550,
		12736	=>	63551,
		12737	=>	63552,
		12738	=>	63553,
		12739	=>	63554,
		12740	=>	63556,
		12741	=>	63557,
		12742	=>	63558,
		12743	=>	63559,
		12744	=>	63560,
		12745	=>	63561,
		12746	=>	63562,
		12747	=>	63563,
		12748	=>	63564,
		12749	=>	63565,
		12750	=>	63566,
		12751	=>	63567,
		12752	=>	63568,
		12753	=>	63569,
		12754	=>	63571,
		12755	=>	63572,
		12756	=>	63573,
		12757	=>	63574,
		12758	=>	63575,
		12759	=>	63576,
		12760	=>	63577,
		12761	=>	63578,
		12762	=>	63579,
		12763	=>	63580,
		12764	=>	63581,
		12765	=>	63582,
		12766	=>	63583,
		12767	=>	63584,
		12768	=>	63586,
		12769	=>	63587,
		12770	=>	63588,
		12771	=>	63589,
		12772	=>	63590,
		12773	=>	63591,
		12774	=>	63592,
		12775	=>	63593,
		12776	=>	63594,
		12777	=>	63595,
		12778	=>	63596,
		12779	=>	63597,
		12780	=>	63598,
		12781	=>	63599,
		12782	=>	63600,
		12783	=>	63602,
		12784	=>	63603,
		12785	=>	63604,
		12786	=>	63605,
		12787	=>	63606,
		12788	=>	63607,
		12789	=>	63608,
		12790	=>	63609,
		12791	=>	63610,
		12792	=>	63611,
		12793	=>	63612,
		12794	=>	63613,
		12795	=>	63614,
		12796	=>	63615,
		12797	=>	63616,
		12798	=>	63617,
		12799	=>	63618,
		12800	=>	63620,
		12801	=>	63621,
		12802	=>	63622,
		12803	=>	63623,
		12804	=>	63624,
		12805	=>	63625,
		12806	=>	63626,
		12807	=>	63627,
		12808	=>	63628,
		12809	=>	63629,
		12810	=>	63630,
		12811	=>	63631,
		12812	=>	63632,
		12813	=>	63633,
		12814	=>	63634,
		12815	=>	63635,
		12816	=>	63636,
		12817	=>	63637,
		12818	=>	63639,
		12819	=>	63640,
		12820	=>	63641,
		12821	=>	63642,
		12822	=>	63643,
		12823	=>	63644,
		12824	=>	63645,
		12825	=>	63646,
		12826	=>	63647,
		12827	=>	63648,
		12828	=>	63649,
		12829	=>	63650,
		12830	=>	63651,
		12831	=>	63652,
		12832	=>	63653,
		12833	=>	63654,
		12834	=>	63655,
		12835	=>	63656,
		12836	=>	63657,
		12837	=>	63659,
		12838	=>	63660,
		12839	=>	63661,
		12840	=>	63662,
		12841	=>	63663,
		12842	=>	63664,
		12843	=>	63665,
		12844	=>	63666,
		12845	=>	63667,
		12846	=>	63668,
		12847	=>	63669,
		12848	=>	63670,
		12849	=>	63671,
		12850	=>	63672,
		12851	=>	63673,
		12852	=>	63674,
		12853	=>	63675,
		12854	=>	63676,
		12855	=>	63677,
		12856	=>	63678,
		12857	=>	63679,
		12858	=>	63680,
		12859	=>	63681,
		12860	=>	63683,
		12861	=>	63684,
		12862	=>	63685,
		12863	=>	63686,
		12864	=>	63687,
		12865	=>	63688,
		12866	=>	63689,
		12867	=>	63690,
		12868	=>	63691,
		12869	=>	63692,
		12870	=>	63693,
		12871	=>	63694,
		12872	=>	63695,
		12873	=>	63696,
		12874	=>	63697,
		12875	=>	63698,
		12876	=>	63699,
		12877	=>	63700,
		12878	=>	63701,
		12879	=>	63702,
		12880	=>	63703,
		12881	=>	63704,
		12882	=>	63705,
		12883	=>	63706,
		12884	=>	63707,
		12885	=>	63708,
		12886	=>	63710,
		12887	=>	63711,
		12888	=>	63712,
		12889	=>	63713,
		12890	=>	63714,
		12891	=>	63715,
		12892	=>	63716,
		12893	=>	63717,
		12894	=>	63718,
		12895	=>	63719,
		12896	=>	63720,
		12897	=>	63721,
		12898	=>	63722,
		12899	=>	63723,
		12900	=>	63724,
		12901	=>	63725,
		12902	=>	63726,
		12903	=>	63727,
		12904	=>	63728,
		12905	=>	63729,
		12906	=>	63730,
		12907	=>	63731,
		12908	=>	63732,
		12909	=>	63733,
		12910	=>	63734,
		12911	=>	63735,
		12912	=>	63736,
		12913	=>	63737,
		12914	=>	63738,
		12915	=>	63739,
		12916	=>	63740,
		12917	=>	63741,
		12918	=>	63742,
		12919	=>	63743,
		12920	=>	63745,
		12921	=>	63746,
		12922	=>	63747,
		12923	=>	63748,
		12924	=>	63749,
		12925	=>	63750,
		12926	=>	63751,
		12927	=>	63752,
		12928	=>	63753,
		12929	=>	63754,
		12930	=>	63755,
		12931	=>	63756,
		12932	=>	63757,
		12933	=>	63758,
		12934	=>	63759,
		12935	=>	63760,
		12936	=>	63761,
		12937	=>	63762,
		12938	=>	63763,
		12939	=>	63764,
		12940	=>	63765,
		12941	=>	63766,
		12942	=>	63767,
		12943	=>	63768,
		12944	=>	63769,
		12945	=>	63770,
		12946	=>	63771,
		12947	=>	63772,
		12948	=>	63773,
		12949	=>	63774,
		12950	=>	63775,
		12951	=>	63776,
		12952	=>	63777,
		12953	=>	63778,
		12954	=>	63779,
		12955	=>	63780,
		12956	=>	63781,
		12957	=>	63782,
		12958	=>	63783,
		12959	=>	63784,
		12960	=>	63785,
		12961	=>	63786,
		12962	=>	63787,
		12963	=>	63788,
		12964	=>	63789,
		12965	=>	63790,
		12966	=>	63791,
		12967	=>	63792,
		12968	=>	63793,
		12969	=>	63794,
		12970	=>	63795,
		12971	=>	63796,
		12972	=>	63797,
		12973	=>	63798,
		12974	=>	63799,
		12975	=>	63800,
		12976	=>	63801,
		12977	=>	63802,
		12978	=>	63803,
		12979	=>	63804,
		12980	=>	63805,
		12981	=>	63806,
		12982	=>	63807,
		12983	=>	63808,
		12984	=>	63809,
		12985	=>	63810,
		12986	=>	63811,
		12987	=>	63812,
		12988	=>	63813,
		12989	=>	63814,
		12990	=>	63816,
		12991	=>	63817,
		12992	=>	63818,
		12993	=>	63819,
		12994	=>	63820,
		12995	=>	63821,
		12996	=>	63822,
		12997	=>	63823,
		12998	=>	63824,
		12999	=>	63825,
		13000	=>	63826,
		13001	=>	63827,
		13002	=>	63828,
		13003	=>	63829,
		13004	=>	63830,
		13005	=>	63831,
		13006	=>	63832,
		13007	=>	63833,
		13008	=>	63834,
		13009	=>	63835,
		13010	=>	63836,
		13011	=>	63837,
		13012	=>	63838,
		13013	=>	63839,
		13014	=>	63840,
		13015	=>	63841,
		13016	=>	63842,
		13017	=>	63843,
		13018	=>	63844,
		13019	=>	63845,
		13020	=>	63846,
		13021	=>	63846,
		13022	=>	63847,
		13023	=>	63848,
		13024	=>	63849,
		13025	=>	63850,
		13026	=>	63851,
		13027	=>	63852,
		13028	=>	63853,
		13029	=>	63854,
		13030	=>	63855,
		13031	=>	63856,
		13032	=>	63857,
		13033	=>	63858,
		13034	=>	63859,
		13035	=>	63860,
		13036	=>	63861,
		13037	=>	63862,
		13038	=>	63863,
		13039	=>	63864,
		13040	=>	63865,
		13041	=>	63866,
		13042	=>	63867,
		13043	=>	63868,
		13044	=>	63869,
		13045	=>	63870,
		13046	=>	63871,
		13047	=>	63872,
		13048	=>	63873,
		13049	=>	63874,
		13050	=>	63875,
		13051	=>	63876,
		13052	=>	63877,
		13053	=>	63878,
		13054	=>	63879,
		13055	=>	63880,
		13056	=>	63881,
		13057	=>	63882,
		13058	=>	63883,
		13059	=>	63884,
		13060	=>	63885,
		13061	=>	63886,
		13062	=>	63887,
		13063	=>	63888,
		13064	=>	63889,
		13065	=>	63890,
		13066	=>	63891,
		13067	=>	63892,
		13068	=>	63893,
		13069	=>	63894,
		13070	=>	63895,
		13071	=>	63896,
		13072	=>	63897,
		13073	=>	63898,
		13074	=>	63899,
		13075	=>	63900,
		13076	=>	63901,
		13077	=>	63902,
		13078	=>	63903,
		13079	=>	63904,
		13080	=>	63905,
		13081	=>	63906,
		13082	=>	63907,
		13083	=>	63908,
		13084	=>	63909,
		13085	=>	63910,
		13086	=>	63911,
		13087	=>	63912,
		13088	=>	63913,
		13089	=>	63914,
		13090	=>	63915,
		13091	=>	63915,
		13092	=>	63916,
		13093	=>	63917,
		13094	=>	63918,
		13095	=>	63919,
		13096	=>	63920,
		13097	=>	63921,
		13098	=>	63922,
		13099	=>	63923,
		13100	=>	63924,
		13101	=>	63925,
		13102	=>	63926,
		13103	=>	63927,
		13104	=>	63928,
		13105	=>	63929,
		13106	=>	63930,
		13107	=>	63931,
		13108	=>	63932,
		13109	=>	63933,
		13110	=>	63934,
		13111	=>	63935,
		13112	=>	63936,
		13113	=>	63937,
		13114	=>	63938,
		13115	=>	63939,
		13116	=>	63940,
		13117	=>	63941,
		13118	=>	63942,
		13119	=>	63943,
		13120	=>	63944,
		13121	=>	63945,
		13122	=>	63946,
		13123	=>	63947,
		13124	=>	63948,
		13125	=>	63948,
		13126	=>	63949,
		13127	=>	63950,
		13128	=>	63951,
		13129	=>	63952,
		13130	=>	63953,
		13131	=>	63954,
		13132	=>	63955,
		13133	=>	63956,
		13134	=>	63957,
		13135	=>	63958,
		13136	=>	63959,
		13137	=>	63960,
		13138	=>	63961,
		13139	=>	63962,
		13140	=>	63963,
		13141	=>	63964,
		13142	=>	63965,
		13143	=>	63966,
		13144	=>	63967,
		13145	=>	63968,
		13146	=>	63969,
		13147	=>	63970,
		13148	=>	63971,
		13149	=>	63972,
		13150	=>	63973,
		13151	=>	63973,
		13152	=>	63974,
		13153	=>	63975,
		13154	=>	63976,
		13155	=>	63977,
		13156	=>	63978,
		13157	=>	63979,
		13158	=>	63980,
		13159	=>	63981,
		13160	=>	63982,
		13161	=>	63983,
		13162	=>	63984,
		13163	=>	63985,
		13164	=>	63986,
		13165	=>	63987,
		13166	=>	63988,
		13167	=>	63989,
		13168	=>	63990,
		13169	=>	63991,
		13170	=>	63992,
		13171	=>	63993,
		13172	=>	63994,
		13173	=>	63995,
		13174	=>	63995,
		13175	=>	63996,
		13176	=>	63997,
		13177	=>	63998,
		13178	=>	63999,
		13179	=>	64000,
		13180	=>	64001,
		13181	=>	64002,
		13182	=>	64003,
		13183	=>	64004,
		13184	=>	64005,
		13185	=>	64006,
		13186	=>	64007,
		13187	=>	64008,
		13188	=>	64009,
		13189	=>	64010,
		13190	=>	64011,
		13191	=>	64012,
		13192	=>	64013,
		13193	=>	64013,
		13194	=>	64014,
		13195	=>	64015,
		13196	=>	64016,
		13197	=>	64017,
		13198	=>	64018,
		13199	=>	64019,
		13200	=>	64020,
		13201	=>	64021,
		13202	=>	64022,
		13203	=>	64023,
		13204	=>	64024,
		13205	=>	64025,
		13206	=>	64026,
		13207	=>	64027,
		13208	=>	64028,
		13209	=>	64029,
		13210	=>	64030,
		13211	=>	64030,
		13212	=>	64031,
		13213	=>	64032,
		13214	=>	64033,
		13215	=>	64034,
		13216	=>	64035,
		13217	=>	64036,
		13218	=>	64037,
		13219	=>	64038,
		13220	=>	64039,
		13221	=>	64040,
		13222	=>	64041,
		13223	=>	64042,
		13224	=>	64043,
		13225	=>	64044,
		13226	=>	64045,
		13227	=>	64045,
		13228	=>	64046,
		13229	=>	64047,
		13230	=>	64048,
		13231	=>	64049,
		13232	=>	64050,
		13233	=>	64051,
		13234	=>	64052,
		13235	=>	64053,
		13236	=>	64054,
		13237	=>	64055,
		13238	=>	64056,
		13239	=>	64057,
		13240	=>	64058,
		13241	=>	64059,
		13242	=>	64060,
		13243	=>	64060,
		13244	=>	64061,
		13245	=>	64062,
		13246	=>	64063,
		13247	=>	64064,
		13248	=>	64065,
		13249	=>	64066,
		13250	=>	64067,
		13251	=>	64068,
		13252	=>	64069,
		13253	=>	64070,
		13254	=>	64071,
		13255	=>	64072,
		13256	=>	64073,
		13257	=>	64073,
		13258	=>	64074,
		13259	=>	64075,
		13260	=>	64076,
		13261	=>	64077,
		13262	=>	64078,
		13263	=>	64079,
		13264	=>	64080,
		13265	=>	64081,
		13266	=>	64082,
		13267	=>	64083,
		13268	=>	64084,
		13269	=>	64085,
		13270	=>	64085,
		13271	=>	64086,
		13272	=>	64087,
		13273	=>	64088,
		13274	=>	64089,
		13275	=>	64090,
		13276	=>	64091,
		13277	=>	64092,
		13278	=>	64093,
		13279	=>	64094,
		13280	=>	64095,
		13281	=>	64096,
		13282	=>	64097,
		13283	=>	64097,
		13284	=>	64098,
		13285	=>	64099,
		13286	=>	64100,
		13287	=>	64101,
		13288	=>	64102,
		13289	=>	64103,
		13290	=>	64104,
		13291	=>	64105,
		13292	=>	64106,
		13293	=>	64107,
		13294	=>	64108,
		13295	=>	64108,
		13296	=>	64109,
		13297	=>	64110,
		13298	=>	64111,
		13299	=>	64112,
		13300	=>	64113,
		13301	=>	64114,
		13302	=>	64115,
		13303	=>	64116,
		13304	=>	64117,
		13305	=>	64118,
		13306	=>	64119,
		13307	=>	64119,
		13308	=>	64120,
		13309	=>	64121,
		13310	=>	64122,
		13311	=>	64123,
		13312	=>	64124,
		13313	=>	64125,
		13314	=>	64126,
		13315	=>	64127,
		13316	=>	64128,
		13317	=>	64129,
		13318	=>	64130,
		13319	=>	64130,
		13320	=>	64131,
		13321	=>	64132,
		13322	=>	64133,
		13323	=>	64134,
		13324	=>	64135,
		13325	=>	64136,
		13326	=>	64137,
		13327	=>	64138,
		13328	=>	64139,
		13329	=>	64140,
		13330	=>	64140,
		13331	=>	64141,
		13332	=>	64142,
		13333	=>	64143,
		13334	=>	64144,
		13335	=>	64145,
		13336	=>	64146,
		13337	=>	64147,
		13338	=>	64148,
		13339	=>	64149,
		13340	=>	64149,
		13341	=>	64150,
		13342	=>	64151,
		13343	=>	64152,
		13344	=>	64153,
		13345	=>	64154,
		13346	=>	64155,
		13347	=>	64156,
		13348	=>	64157,
		13349	=>	64158,
		13350	=>	64158,
		13351	=>	64159,
		13352	=>	64160,
		13353	=>	64161,
		13354	=>	64162,
		13355	=>	64163,
		13356	=>	64164,
		13357	=>	64165,
		13358	=>	64166,
		13359	=>	64167,
		13360	=>	64167,
		13361	=>	64168,
		13362	=>	64169,
		13363	=>	64170,
		13364	=>	64171,
		13365	=>	64172,
		13366	=>	64173,
		13367	=>	64174,
		13368	=>	64175,
		13369	=>	64176,
		13370	=>	64176,
		13371	=>	64177,
		13372	=>	64178,
		13373	=>	64179,
		13374	=>	64180,
		13375	=>	64181,
		13376	=>	64182,
		13377	=>	64183,
		13378	=>	64184,
		13379	=>	64184,
		13380	=>	64185,
		13381	=>	64186,
		13382	=>	64187,
		13383	=>	64188,
		13384	=>	64189,
		13385	=>	64190,
		13386	=>	64191,
		13387	=>	64192,
		13388	=>	64193,
		13389	=>	64193,
		13390	=>	64194,
		13391	=>	64195,
		13392	=>	64196,
		13393	=>	64197,
		13394	=>	64198,
		13395	=>	64199,
		13396	=>	64200,
		13397	=>	64201,
		13398	=>	64201,
		13399	=>	64202,
		13400	=>	64203,
		13401	=>	64204,
		13402	=>	64205,
		13403	=>	64206,
		13404	=>	64207,
		13405	=>	64208,
		13406	=>	64208,
		13407	=>	64209,
		13408	=>	64210,
		13409	=>	64211,
		13410	=>	64212,
		13411	=>	64213,
		13412	=>	64214,
		13413	=>	64215,
		13414	=>	64216,
		13415	=>	64216,
		13416	=>	64217,
		13417	=>	64218,
		13418	=>	64219,
		13419	=>	64220,
		13420	=>	64221,
		13421	=>	64222,
		13422	=>	64223,
		13423	=>	64223,
		13424	=>	64224,
		13425	=>	64225,
		13426	=>	64226,
		13427	=>	64227,
		13428	=>	64228,
		13429	=>	64229,
		13430	=>	64230,
		13431	=>	64231,
		13432	=>	64231,
		13433	=>	64232,
		13434	=>	64233,
		13435	=>	64234,
		13436	=>	64235,
		13437	=>	64236,
		13438	=>	64237,
		13439	=>	64238,
		13440	=>	64238,
		13441	=>	64239,
		13442	=>	64240,
		13443	=>	64241,
		13444	=>	64242,
		13445	=>	64243,
		13446	=>	64244,
		13447	=>	64245,
		13448	=>	64245,
		13449	=>	64246,
		13450	=>	64247,
		13451	=>	64248,
		13452	=>	64249,
		13453	=>	64250,
		13454	=>	64251,
		13455	=>	64251,
		13456	=>	64252,
		13457	=>	64253,
		13458	=>	64254,
		13459	=>	64255,
		13460	=>	64256,
		13461	=>	64257,
		13462	=>	64258,
		13463	=>	64258,
		13464	=>	64259,
		13465	=>	64260,
		13466	=>	64261,
		13467	=>	64262,
		13468	=>	64263,
		13469	=>	64264,
		13470	=>	64265,
		13471	=>	64265,
		13472	=>	64266,
		13473	=>	64267,
		13474	=>	64268,
		13475	=>	64269,
		13476	=>	64270,
		13477	=>	64271,
		13478	=>	64271,
		13479	=>	64272,
		13480	=>	64273,
		13481	=>	64274,
		13482	=>	64275,
		13483	=>	64276,
		13484	=>	64277,
		13485	=>	64277,
		13486	=>	64278,
		13487	=>	64279,
		13488	=>	64280,
		13489	=>	64281,
		13490	=>	64282,
		13491	=>	64283,
		13492	=>	64284,
		13493	=>	64284,
		13494	=>	64285,
		13495	=>	64286,
		13496	=>	64287,
		13497	=>	64288,
		13498	=>	64289,
		13499	=>	64290,
		13500	=>	64290,
		13501	=>	64291,
		13502	=>	64292,
		13503	=>	64293,
		13504	=>	64294,
		13505	=>	64295,
		13506	=>	64296,
		13507	=>	64296,
		13508	=>	64297,
		13509	=>	64298,
		13510	=>	64299,
		13511	=>	64300,
		13512	=>	64301,
		13513	=>	64302,
		13514	=>	64302,
		13515	=>	64303,
		13516	=>	64304,
		13517	=>	64305,
		13518	=>	64306,
		13519	=>	64307,
		13520	=>	64307,
		13521	=>	64308,
		13522	=>	64309,
		13523	=>	64310,
		13524	=>	64311,
		13525	=>	64312,
		13526	=>	64313,
		13527	=>	64313,
		13528	=>	64314,
		13529	=>	64315,
		13530	=>	64316,
		13531	=>	64317,
		13532	=>	64318,
		13533	=>	64319,
		13534	=>	64319,
		13535	=>	64320,
		13536	=>	64321,
		13537	=>	64322,
		13538	=>	64323,
		13539	=>	64324,
		13540	=>	64324,
		13541	=>	64325,
		13542	=>	64326,
		13543	=>	64327,
		13544	=>	64328,
		13545	=>	64329,
		13546	=>	64330,
		13547	=>	64330,
		13548	=>	64331,
		13549	=>	64332,
		13550	=>	64333,
		13551	=>	64334,
		13552	=>	64335,
		13553	=>	64335,
		13554	=>	64336,
		13555	=>	64337,
		13556	=>	64338,
		13557	=>	64339,
		13558	=>	64340,
		13559	=>	64340,
		13560	=>	64341,
		13561	=>	64342,
		13562	=>	64343,
		13563	=>	64344,
		13564	=>	64345,
		13565	=>	64346,
		13566	=>	64346,
		13567	=>	64347,
		13568	=>	64348,
		13569	=>	64349,
		13570	=>	64350,
		13571	=>	64351,
		13572	=>	64351,
		13573	=>	64352,
		13574	=>	64353,
		13575	=>	64354,
		13576	=>	64355,
		13577	=>	64356,
		13578	=>	64356,
		13579	=>	64357,
		13580	=>	64358,
		13581	=>	64359,
		13582	=>	64360,
		13583	=>	64361,
		13584	=>	64361,
		13585	=>	64362,
		13586	=>	64363,
		13587	=>	64364,
		13588	=>	64365,
		13589	=>	64366,
		13590	=>	64366,
		13591	=>	64367,
		13592	=>	64368,
		13593	=>	64369,
		13594	=>	64370,
		13595	=>	64371,
		13596	=>	64371,
		13597	=>	64372,
		13598	=>	64373,
		13599	=>	64374,
		13600	=>	64375,
		13601	=>	64376,
		13602	=>	64376,
		13603	=>	64377,
		13604	=>	64378,
		13605	=>	64379,
		13606	=>	64380,
		13607	=>	64380,
		13608	=>	64381,
		13609	=>	64382,
		13610	=>	64383,
		13611	=>	64384,
		13612	=>	64385,
		13613	=>	64385,
		13614	=>	64386,
		13615	=>	64387,
		13616	=>	64388,
		13617	=>	64389,
		13618	=>	64390,
		13619	=>	64390,
		13620	=>	64391,
		13621	=>	64392,
		13622	=>	64393,
		13623	=>	64394,
		13624	=>	64394,
		13625	=>	64395,
		13626	=>	64396,
		13627	=>	64397,
		13628	=>	64398,
		13629	=>	64399,
		13630	=>	64399,
		13631	=>	64400,
		13632	=>	64401,
		13633	=>	64402,
		13634	=>	64403,
		13635	=>	64404,
		13636	=>	64404,
		13637	=>	64405,
		13638	=>	64406,
		13639	=>	64407,
		13640	=>	64408,
		13641	=>	64408,
		13642	=>	64409,
		13643	=>	64410,
		13644	=>	64411,
		13645	=>	64412,
		13646	=>	64413,
		13647	=>	64413,
		13648	=>	64414,
		13649	=>	64415,
		13650	=>	64416,
		13651	=>	64417,
		13652	=>	64417,
		13653	=>	64418,
		13654	=>	64419,
		13655	=>	64420,
		13656	=>	64421,
		13657	=>	64421,
		13658	=>	64422,
		13659	=>	64423,
		13660	=>	64424,
		13661	=>	64425,
		13662	=>	64426,
		13663	=>	64426,
		13664	=>	64427,
		13665	=>	64428,
		13666	=>	64429,
		13667	=>	64430,
		13668	=>	64430,
		13669	=>	64431,
		13670	=>	64432,
		13671	=>	64433,
		13672	=>	64434,
		13673	=>	64434,
		13674	=>	64435,
		13675	=>	64436,
		13676	=>	64437,
		13677	=>	64438,
		13678	=>	64438,
		13679	=>	64439,
		13680	=>	64440,
		13681	=>	64441,
		13682	=>	64442,
		13683	=>	64442,
		13684	=>	64443,
		13685	=>	64444,
		13686	=>	64445,
		13687	=>	64446,
		13688	=>	64446,
		13689	=>	64447,
		13690	=>	64448,
		13691	=>	64449,
		13692	=>	64450,
		13693	=>	64450,
		13694	=>	64451,
		13695	=>	64452,
		13696	=>	64453,
		13697	=>	64454,
		13698	=>	64455,
		13699	=>	64455,
		13700	=>	64456,
		13701	=>	64457,
		13702	=>	64458,
		13703	=>	64458,
		13704	=>	64459,
		13705	=>	64460,
		13706	=>	64461,
		13707	=>	64462,
		13708	=>	64462,
		13709	=>	64463,
		13710	=>	64464,
		13711	=>	64465,
		13712	=>	64466,
		13713	=>	64466,
		13714	=>	64467,
		13715	=>	64468,
		13716	=>	64469,
		13717	=>	64470,
		13718	=>	64470,
		13719	=>	64471,
		13720	=>	64472,
		13721	=>	64473,
		13722	=>	64474,
		13723	=>	64474,
		13724	=>	64475,
		13725	=>	64476,
		13726	=>	64477,
		13727	=>	64478,
		13728	=>	64478,
		13729	=>	64479,
		13730	=>	64480,
		13731	=>	64481,
		13732	=>	64482,
		13733	=>	64482,
		13734	=>	64483,
		13735	=>	64484,
		13736	=>	64485,
		13737	=>	64485,
		13738	=>	64486,
		13739	=>	64487,
		13740	=>	64488,
		13741	=>	64489,
		13742	=>	64489,
		13743	=>	64490,
		13744	=>	64491,
		13745	=>	64492,
		13746	=>	64493,
		13747	=>	64493,
		13748	=>	64494,
		13749	=>	64495,
		13750	=>	64496,
		13751	=>	64496,
		13752	=>	64497,
		13753	=>	64498,
		13754	=>	64499,
		13755	=>	64500,
		13756	=>	64500,
		13757	=>	64501,
		13758	=>	64502,
		13759	=>	64503,
		13760	=>	64504,
		13761	=>	64504,
		13762	=>	64505,
		13763	=>	64506,
		13764	=>	64507,
		13765	=>	64507,
		13766	=>	64508,
		13767	=>	64509,
		13768	=>	64510,
		13769	=>	64511,
		13770	=>	64511,
		13771	=>	64512,
		13772	=>	64513,
		13773	=>	64514,
		13774	=>	64514,
		13775	=>	64515,
		13776	=>	64516,
		13777	=>	64517,
		13778	=>	64518,
		13779	=>	64518,
		13780	=>	64519,
		13781	=>	64520,
		13782	=>	64521,
		13783	=>	64521,
		13784	=>	64522,
		13785	=>	64523,
		13786	=>	64524,
		13787	=>	64525,
		13788	=>	64525,
		13789	=>	64526,
		13790	=>	64527,
		13791	=>	64528,
		13792	=>	64528,
		13793	=>	64529,
		13794	=>	64530,
		13795	=>	64531,
		13796	=>	64532,
		13797	=>	64532,
		13798	=>	64533,
		13799	=>	64534,
		13800	=>	64535,
		13801	=>	64535,
		13802	=>	64536,
		13803	=>	64537,
		13804	=>	64538,
		13805	=>	64538,
		13806	=>	64539,
		13807	=>	64540,
		13808	=>	64541,
		13809	=>	64542,
		13810	=>	64542,
		13811	=>	64543,
		13812	=>	64544,
		13813	=>	64545,
		13814	=>	64545,
		13815	=>	64546,
		13816	=>	64547,
		13817	=>	64548,
		13818	=>	64548,
		13819	=>	64549,
		13820	=>	64550,
		13821	=>	64551,
		13822	=>	64551,
		13823	=>	64552,
		13824	=>	64553,
		13825	=>	64554,
		13826	=>	64555,
		13827	=>	64555,
		13828	=>	64556,
		13829	=>	64557,
		13830	=>	64558,
		13831	=>	64558,
		13832	=>	64559,
		13833	=>	64560,
		13834	=>	64561,
		13835	=>	64561,
		13836	=>	64562,
		13837	=>	64563,
		13838	=>	64564,
		13839	=>	64564,
		13840	=>	64565,
		13841	=>	64566,
		13842	=>	64567,
		13843	=>	64567,
		13844	=>	64568,
		13845	=>	64569,
		13846	=>	64570,
		13847	=>	64570,
		13848	=>	64571,
		13849	=>	64572,
		13850	=>	64573,
		13851	=>	64574,
		13852	=>	64574,
		13853	=>	64575,
		13854	=>	64576,
		13855	=>	64577,
		13856	=>	64577,
		13857	=>	64578,
		13858	=>	64579,
		13859	=>	64580,
		13860	=>	64580,
		13861	=>	64581,
		13862	=>	64582,
		13863	=>	64583,
		13864	=>	64583,
		13865	=>	64584,
		13866	=>	64585,
		13867	=>	64586,
		13868	=>	64586,
		13869	=>	64587,
		13870	=>	64588,
		13871	=>	64589,
		13872	=>	64589,
		13873	=>	64590,
		13874	=>	64591,
		13875	=>	64592,
		13876	=>	64592,
		13877	=>	64593,
		13878	=>	64594,
		13879	=>	64595,
		13880	=>	64595,
		13881	=>	64596,
		13882	=>	64597,
		13883	=>	64598,
		13884	=>	64598,
		13885	=>	64599,
		13886	=>	64600,
		13887	=>	64601,
		13888	=>	64601,
		13889	=>	64602,
		13890	=>	64603,
		13891	=>	64603,
		13892	=>	64604,
		13893	=>	64605,
		13894	=>	64606,
		13895	=>	64606,
		13896	=>	64607,
		13897	=>	64608,
		13898	=>	64609,
		13899	=>	64609,
		13900	=>	64610,
		13901	=>	64611,
		13902	=>	64612,
		13903	=>	64612,
		13904	=>	64613,
		13905	=>	64614,
		13906	=>	64615,
		13907	=>	64615,
		13908	=>	64616,
		13909	=>	64617,
		13910	=>	64618,
		13911	=>	64618,
		13912	=>	64619,
		13913	=>	64620,
		13914	=>	64621,
		13915	=>	64621,
		13916	=>	64622,
		13917	=>	64623,
		13918	=>	64623,
		13919	=>	64624,
		13920	=>	64625,
		13921	=>	64626,
		13922	=>	64626,
		13923	=>	64627,
		13924	=>	64628,
		13925	=>	64629,
		13926	=>	64629,
		13927	=>	64630,
		13928	=>	64631,
		13929	=>	64632,
		13930	=>	64632,
		13931	=>	64633,
		13932	=>	64634,
		13933	=>	64634,
		13934	=>	64635,
		13935	=>	64636,
		13936	=>	64637,
		13937	=>	64637,
		13938	=>	64638,
		13939	=>	64639,
		13940	=>	64640,
		13941	=>	64640,
		13942	=>	64641,
		13943	=>	64642,
		13944	=>	64642,
		13945	=>	64643,
		13946	=>	64644,
		13947	=>	64645,
		13948	=>	64645,
		13949	=>	64646,
		13950	=>	64647,
		13951	=>	64648,
		13952	=>	64648,
		13953	=>	64649,
		13954	=>	64650,
		13955	=>	64650,
		13956	=>	64651,
		13957	=>	64652,
		13958	=>	64653,
		13959	=>	64653,
		13960	=>	64654,
		13961	=>	64655,
		13962	=>	64656,
		13963	=>	64656,
		13964	=>	64657,
		13965	=>	64658,
		13966	=>	64658,
		13967	=>	64659,
		13968	=>	64660,
		13969	=>	64661,
		13970	=>	64661,
		13971	=>	64662,
		13972	=>	64663,
		13973	=>	64663,
		13974	=>	64664,
		13975	=>	64665,
		13976	=>	64666,
		13977	=>	64666,
		13978	=>	64667,
		13979	=>	64668,
		13980	=>	64669,
		13981	=>	64669,
		13982	=>	64670,
		13983	=>	64671,
		13984	=>	64671,
		13985	=>	64672,
		13986	=>	64673,
		13987	=>	64674,
		13988	=>	64674,
		13989	=>	64675,
		13990	=>	64676,
		13991	=>	64676,
		13992	=>	64677,
		13993	=>	64678,
		13994	=>	64679,
		13995	=>	64679,
		13996	=>	64680,
		13997	=>	64681,
		13998	=>	64681,
		13999	=>	64682,
		14000	=>	64683,
		14001	=>	64684,
		14002	=>	64684,
		14003	=>	64685,
		14004	=>	64686,
		14005	=>	64686,
		14006	=>	64687,
		14007	=>	64688,
		14008	=>	64688,
		14009	=>	64689,
		14010	=>	64690,
		14011	=>	64691,
		14012	=>	64691,
		14013	=>	64692,
		14014	=>	64693,
		14015	=>	64693,
		14016	=>	64694,
		14017	=>	64695,
		14018	=>	64696,
		14019	=>	64696,
		14020	=>	64697,
		14021	=>	64698,
		14022	=>	64698,
		14023	=>	64699,
		14024	=>	64700,
		14025	=>	64701,
		14026	=>	64701,
		14027	=>	64702,
		14028	=>	64703,
		14029	=>	64703,
		14030	=>	64704,
		14031	=>	64705,
		14032	=>	64705,
		14033	=>	64706,
		14034	=>	64707,
		14035	=>	64708,
		14036	=>	64708,
		14037	=>	64709,
		14038	=>	64710,
		14039	=>	64710,
		14040	=>	64711,
		14041	=>	64712,
		14042	=>	64712,
		14043	=>	64713,
		14044	=>	64714,
		14045	=>	64715,
		14046	=>	64715,
		14047	=>	64716,
		14048	=>	64717,
		14049	=>	64717,
		14050	=>	64718,
		14051	=>	64719,
		14052	=>	64719,
		14053	=>	64720,
		14054	=>	64721,
		14055	=>	64722,
		14056	=>	64722,
		14057	=>	64723,
		14058	=>	64724,
		14059	=>	64724,
		14060	=>	64725,
		14061	=>	64726,
		14062	=>	64726,
		14063	=>	64727,
		14064	=>	64728,
		14065	=>	64728,
		14066	=>	64729,
		14067	=>	64730,
		14068	=>	64731,
		14069	=>	64731,
		14070	=>	64732,
		14071	=>	64733,
		14072	=>	64733,
		14073	=>	64734,
		14074	=>	64735,
		14075	=>	64735,
		14076	=>	64736,
		14077	=>	64737,
		14078	=>	64737,
		14079	=>	64738,
		14080	=>	64739,
		14081	=>	64740,
		14082	=>	64740,
		14083	=>	64741,
		14084	=>	64742,
		14085	=>	64742,
		14086	=>	64743,
		14087	=>	64744,
		14088	=>	64744,
		14089	=>	64745,
		14090	=>	64746,
		14091	=>	64746,
		14092	=>	64747,
		14093	=>	64748,
		14094	=>	64748,
		14095	=>	64749,
		14096	=>	64750,
		14097	=>	64750,
		14098	=>	64751,
		14099	=>	64752,
		14100	=>	64753,
		14101	=>	64753,
		14102	=>	64754,
		14103	=>	64755,
		14104	=>	64755,
		14105	=>	64756,
		14106	=>	64757,
		14107	=>	64757,
		14108	=>	64758,
		14109	=>	64759,
		14110	=>	64759,
		14111	=>	64760,
		14112	=>	64761,
		14113	=>	64761,
		14114	=>	64762,
		14115	=>	64763,
		14116	=>	64763,
		14117	=>	64764,
		14118	=>	64765,
		14119	=>	64765,
		14120	=>	64766,
		14121	=>	64767,
		14122	=>	64767,
		14123	=>	64768,
		14124	=>	64769,
		14125	=>	64769,
		14126	=>	64770,
		14127	=>	64771,
		14128	=>	64772,
		14129	=>	64772,
		14130	=>	64773,
		14131	=>	64774,
		14132	=>	64774,
		14133	=>	64775,
		14134	=>	64776,
		14135	=>	64776,
		14136	=>	64777,
		14137	=>	64778,
		14138	=>	64778,
		14139	=>	64779,
		14140	=>	64780,
		14141	=>	64780,
		14142	=>	64781,
		14143	=>	64782,
		14144	=>	64782,
		14145	=>	64783,
		14146	=>	64784,
		14147	=>	64784,
		14148	=>	64785,
		14149	=>	64786,
		14150	=>	64786,
		14151	=>	64787,
		14152	=>	64788,
		14153	=>	64788,
		14154	=>	64789,
		14155	=>	64790,
		14156	=>	64790,
		14157	=>	64791,
		14158	=>	64792,
		14159	=>	64792,
		14160	=>	64793,
		14161	=>	64794,
		14162	=>	64794,
		14163	=>	64795,
		14164	=>	64796,
		14165	=>	64796,
		14166	=>	64797,
		14167	=>	64798,
		14168	=>	64798,
		14169	=>	64799,
		14170	=>	64800,
		14171	=>	64800,
		14172	=>	64801,
		14173	=>	64802,
		14174	=>	64802,
		14175	=>	64803,
		14176	=>	64804,
		14177	=>	64804,
		14178	=>	64805,
		14179	=>	64806,
		14180	=>	64806,
		14181	=>	64807,
		14182	=>	64807,
		14183	=>	64808,
		14184	=>	64809,
		14185	=>	64809,
		14186	=>	64810,
		14187	=>	64811,
		14188	=>	64811,
		14189	=>	64812,
		14190	=>	64813,
		14191	=>	64813,
		14192	=>	64814,
		14193	=>	64815,
		14194	=>	64815,
		14195	=>	64816,
		14196	=>	64817,
		14197	=>	64817,
		14198	=>	64818,
		14199	=>	64819,
		14200	=>	64819,
		14201	=>	64820,
		14202	=>	64821,
		14203	=>	64821,
		14204	=>	64822,
		14205	=>	64823,
		14206	=>	64823,
		14207	=>	64824,
		14208	=>	64825,
		14209	=>	64825,
		14210	=>	64826,
		14211	=>	64826,
		14212	=>	64827,
		14213	=>	64828,
		14214	=>	64828,
		14215	=>	64829,
		14216	=>	64830,
		14217	=>	64830,
		14218	=>	64831,
		14219	=>	64832,
		14220	=>	64832,
		14221	=>	64833,
		14222	=>	64834,
		14223	=>	64834,
		14224	=>	64835,
		14225	=>	64836,
		14226	=>	64836,
		14227	=>	64837,
		14228	=>	64837,
		14229	=>	64838,
		14230	=>	64839,
		14231	=>	64839,
		14232	=>	64840,
		14233	=>	64841,
		14234	=>	64841,
		14235	=>	64842,
		14236	=>	64843,
		14237	=>	64843,
		14238	=>	64844,
		14239	=>	64845,
		14240	=>	64845,
		14241	=>	64846,
		14242	=>	64846,
		14243	=>	64847,
		14244	=>	64848,
		14245	=>	64848,
		14246	=>	64849,
		14247	=>	64850,
		14248	=>	64850,
		14249	=>	64851,
		14250	=>	64852,
		14251	=>	64852,
		14252	=>	64853,
		14253	=>	64853,
		14254	=>	64854,
		14255	=>	64855,
		14256	=>	64855,
		14257	=>	64856,
		14258	=>	64857,
		14259	=>	64857,
		14260	=>	64858,
		14261	=>	64859,
		14262	=>	64859,
		14263	=>	64860,
		14264	=>	64860,
		14265	=>	64861,
		14266	=>	64862,
		14267	=>	64862,
		14268	=>	64863,
		14269	=>	64864,
		14270	=>	64864,
		14271	=>	64865,
		14272	=>	64866,
		14273	=>	64866,
		14274	=>	64867,
		14275	=>	64867,
		14276	=>	64868,
		14277	=>	64869,
		14278	=>	64869,
		14279	=>	64870,
		14280	=>	64871,
		14281	=>	64871,
		14282	=>	64872,
		14283	=>	64872,
		14284	=>	64873,
		14285	=>	64874,
		14286	=>	64874,
		14287	=>	64875,
		14288	=>	64876,
		14289	=>	64876,
		14290	=>	64877,
		14291	=>	64878,
		14292	=>	64878,
		14293	=>	64879,
		14294	=>	64879,
		14295	=>	64880,
		14296	=>	64881,
		14297	=>	64881,
		14298	=>	64882,
		14299	=>	64883,
		14300	=>	64883,
		14301	=>	64884,
		14302	=>	64884,
		14303	=>	64885,
		14304	=>	64886,
		14305	=>	64886,
		14306	=>	64887,
		14307	=>	64887,
		14308	=>	64888,
		14309	=>	64889,
		14310	=>	64889,
		14311	=>	64890,
		14312	=>	64891,
		14313	=>	64891,
		14314	=>	64892,
		14315	=>	64892,
		14316	=>	64893,
		14317	=>	64894,
		14318	=>	64894,
		14319	=>	64895,
		14320	=>	64896,
		14321	=>	64896,
		14322	=>	64897,
		14323	=>	64897,
		14324	=>	64898,
		14325	=>	64899,
		14326	=>	64899,
		14327	=>	64900,
		14328	=>	64900,
		14329	=>	64901,
		14330	=>	64902,
		14331	=>	64902,
		14332	=>	64903,
		14333	=>	64904,
		14334	=>	64904,
		14335	=>	64905,
		14336	=>	64905,
		14337	=>	64906,
		14338	=>	64907,
		14339	=>	64907,
		14340	=>	64908,
		14341	=>	64908,
		14342	=>	64909,
		14343	=>	64910,
		14344	=>	64910,
		14345	=>	64911,
		14346	=>	64911,
		14347	=>	64912,
		14348	=>	64913,
		14349	=>	64913,
		14350	=>	64914,
		14351	=>	64915,
		14352	=>	64915,
		14353	=>	64916,
		14354	=>	64916,
		14355	=>	64917,
		14356	=>	64918,
		14357	=>	64918,
		14358	=>	64919,
		14359	=>	64919,
		14360	=>	64920,
		14361	=>	64921,
		14362	=>	64921,
		14363	=>	64922,
		14364	=>	64922,
		14365	=>	64923,
		14366	=>	64924,
		14367	=>	64924,
		14368	=>	64925,
		14369	=>	64925,
		14370	=>	64926,
		14371	=>	64927,
		14372	=>	64927,
		14373	=>	64928,
		14374	=>	64928,
		14375	=>	64929,
		14376	=>	64930,
		14377	=>	64930,
		14378	=>	64931,
		14379	=>	64931,
		14380	=>	64932,
		14381	=>	64933,
		14382	=>	64933,
		14383	=>	64934,
		14384	=>	64934,
		14385	=>	64935,
		14386	=>	64936,
		14387	=>	64936,
		14388	=>	64937,
		14389	=>	64937,
		14390	=>	64938,
		14391	=>	64939,
		14392	=>	64939,
		14393	=>	64940,
		14394	=>	64940,
		14395	=>	64941,
		14396	=>	64942,
		14397	=>	64942,
		14398	=>	64943,
		14399	=>	64943,
		14400	=>	64944,
		14401	=>	64945,
		14402	=>	64945,
		14403	=>	64946,
		14404	=>	64946,
		14405	=>	64947,
		14406	=>	64948,
		14407	=>	64948,
		14408	=>	64949,
		14409	=>	64949,
		14410	=>	64950,
		14411	=>	64951,
		14412	=>	64951,
		14413	=>	64952,
		14414	=>	64952,
		14415	=>	64953,
		14416	=>	64953,
		14417	=>	64954,
		14418	=>	64955,
		14419	=>	64955,
		14420	=>	64956,
		14421	=>	64956,
		14422	=>	64957,
		14423	=>	64958,
		14424	=>	64958,
		14425	=>	64959,
		14426	=>	64959,
		14427	=>	64960,
		14428	=>	64961,
		14429	=>	64961,
		14430	=>	64962,
		14431	=>	64962,
		14432	=>	64963,
		14433	=>	64963,
		14434	=>	64964,
		14435	=>	64965,
		14436	=>	64965,
		14437	=>	64966,
		14438	=>	64966,
		14439	=>	64967,
		14440	=>	64968,
		14441	=>	64968,
		14442	=>	64969,
		14443	=>	64969,
		14444	=>	64970,
		14445	=>	64970,
		14446	=>	64971,
		14447	=>	64972,
		14448	=>	64972,
		14449	=>	64973,
		14450	=>	64973,
		14451	=>	64974,
		14452	=>	64974,
		14453	=>	64975,
		14454	=>	64976,
		14455	=>	64976,
		14456	=>	64977,
		14457	=>	64977,
		14458	=>	64978,
		14459	=>	64979,
		14460	=>	64979,
		14461	=>	64980,
		14462	=>	64980,
		14463	=>	64981,
		14464	=>	64981,
		14465	=>	64982,
		14466	=>	64983,
		14467	=>	64983,
		14468	=>	64984,
		14469	=>	64984,
		14470	=>	64985,
		14471	=>	64985,
		14472	=>	64986,
		14473	=>	64987,
		14474	=>	64987,
		14475	=>	64988,
		14476	=>	64988,
		14477	=>	64989,
		14478	=>	64989,
		14479	=>	64990,
		14480	=>	64991,
		14481	=>	64991,
		14482	=>	64992,
		14483	=>	64992,
		14484	=>	64993,
		14485	=>	64993,
		14486	=>	64994,
		14487	=>	64995,
		14488	=>	64995,
		14489	=>	64996,
		14490	=>	64996,
		14491	=>	64997,
		14492	=>	64997,
		14493	=>	64998,
		14494	=>	64999,
		14495	=>	64999,
		14496	=>	65000,
		14497	=>	65000,
		14498	=>	65001,
		14499	=>	65001,
		14500	=>	65002,
		14501	=>	65002,
		14502	=>	65003,
		14503	=>	65004,
		14504	=>	65004,
		14505	=>	65005,
		14506	=>	65005,
		14507	=>	65006,
		14508	=>	65006,
		14509	=>	65007,
		14510	=>	65008,
		14511	=>	65008,
		14512	=>	65009,
		14513	=>	65009,
		14514	=>	65010,
		14515	=>	65010,
		14516	=>	65011,
		14517	=>	65011,
		14518	=>	65012,
		14519	=>	65013,
		14520	=>	65013,
		14521	=>	65014,
		14522	=>	65014,
		14523	=>	65015,
		14524	=>	65015,
		14525	=>	65016,
		14526	=>	65016,
		14527	=>	65017,
		14528	=>	65018,
		14529	=>	65018,
		14530	=>	65019,
		14531	=>	65019,
		14532	=>	65020,
		14533	=>	65020,
		14534	=>	65021,
		14535	=>	65021,
		14536	=>	65022,
		14537	=>	65023,
		14538	=>	65023,
		14539	=>	65024,
		14540	=>	65024,
		14541	=>	65025,
		14542	=>	65025,
		14543	=>	65026,
		14544	=>	65026,
		14545	=>	65027,
		14546	=>	65028,
		14547	=>	65028,
		14548	=>	65029,
		14549	=>	65029,
		14550	=>	65030,
		14551	=>	65030,
		14552	=>	65031,
		14553	=>	65031,
		14554	=>	65032,
		14555	=>	65033,
		14556	=>	65033,
		14557	=>	65034,
		14558	=>	65034,
		14559	=>	65035,
		14560	=>	65035,
		14561	=>	65036,
		14562	=>	65036,
		14563	=>	65037,
		14564	=>	65037,
		14565	=>	65038,
		14566	=>	65039,
		14567	=>	65039,
		14568	=>	65040,
		14569	=>	65040,
		14570	=>	65041,
		14571	=>	65041,
		14572	=>	65042,
		14573	=>	65042,
		14574	=>	65043,
		14575	=>	65043,
		14576	=>	65044,
		14577	=>	65044,
		14578	=>	65045,
		14579	=>	65046,
		14580	=>	65046,
		14581	=>	65047,
		14582	=>	65047,
		14583	=>	65048,
		14584	=>	65048,
		14585	=>	65049,
		14586	=>	65049,
		14587	=>	65050,
		14588	=>	65050,
		14589	=>	65051,
		14590	=>	65052,
		14591	=>	65052,
		14592	=>	65053,
		14593	=>	65053,
		14594	=>	65054,
		14595	=>	65054,
		14596	=>	65055,
		14597	=>	65055,
		14598	=>	65056,
		14599	=>	65056,
		14600	=>	65057,
		14601	=>	65057,
		14602	=>	65058,
		14603	=>	65058,
		14604	=>	65059,
		14605	=>	65060,
		14606	=>	65060,
		14607	=>	65061,
		14608	=>	65061,
		14609	=>	65062,
		14610	=>	65062,
		14611	=>	65063,
		14612	=>	65063,
		14613	=>	65064,
		14614	=>	65064,
		14615	=>	65065,
		14616	=>	65065,
		14617	=>	65066,
		14618	=>	65066,
		14619	=>	65067,
		14620	=>	65068,
		14621	=>	65068,
		14622	=>	65069,
		14623	=>	65069,
		14624	=>	65070,
		14625	=>	65070,
		14626	=>	65071,
		14627	=>	65071,
		14628	=>	65072,
		14629	=>	65072,
		14630	=>	65073,
		14631	=>	65073,
		14632	=>	65074,
		14633	=>	65074,
		14634	=>	65075,
		14635	=>	65075,
		14636	=>	65076,
		14637	=>	65076,
		14638	=>	65077,
		14639	=>	65078,
		14640	=>	65078,
		14641	=>	65079,
		14642	=>	65079,
		14643	=>	65080,
		14644	=>	65080,
		14645	=>	65081,
		14646	=>	65081,
		14647	=>	65082,
		14648	=>	65082,
		14649	=>	65083,
		14650	=>	65083,
		14651	=>	65084,
		14652	=>	65084,
		14653	=>	65085,
		14654	=>	65085,
		14655	=>	65086,
		14656	=>	65086,
		14657	=>	65087,
		14658	=>	65087,
		14659	=>	65088,
		14660	=>	65088,
		14661	=>	65089,
		14662	=>	65089,
		14663	=>	65090,
		14664	=>	65090,
		14665	=>	65091,
		14666	=>	65092,
		14667	=>	65092,
		14668	=>	65093,
		14669	=>	65093,
		14670	=>	65094,
		14671	=>	65094,
		14672	=>	65095,
		14673	=>	65095,
		14674	=>	65096,
		14675	=>	65096,
		14676	=>	65097,
		14677	=>	65097,
		14678	=>	65098,
		14679	=>	65098,
		14680	=>	65099,
		14681	=>	65099,
		14682	=>	65100,
		14683	=>	65100,
		14684	=>	65101,
		14685	=>	65101,
		14686	=>	65102,
		14687	=>	65102,
		14688	=>	65103,
		14689	=>	65103,
		14690	=>	65104,
		14691	=>	65104,
		14692	=>	65105,
		14693	=>	65105,
		14694	=>	65106,
		14695	=>	65106,
		14696	=>	65107,
		14697	=>	65107,
		14698	=>	65108,
		14699	=>	65108,
		14700	=>	65109,
		14701	=>	65109,
		14702	=>	65110,
		14703	=>	65110,
		14704	=>	65111,
		14705	=>	65111,
		14706	=>	65112,
		14707	=>	65112,
		14708	=>	65113,
		14709	=>	65113,
		14710	=>	65114,
		14711	=>	65114,
		14712	=>	65115,
		14713	=>	65115,
		14714	=>	65116,
		14715	=>	65116,
		14716	=>	65117,
		14717	=>	65117,
		14718	=>	65118,
		14719	=>	65118,
		14720	=>	65119,
		14721	=>	65119,
		14722	=>	65120,
		14723	=>	65120,
		14724	=>	65121,
		14725	=>	65121,
		14726	=>	65122,
		14727	=>	65122,
		14728	=>	65123,
		14729	=>	65123,
		14730	=>	65124,
		14731	=>	65124,
		14732	=>	65125,
		14733	=>	65125,
		14734	=>	65126,
		14735	=>	65126,
		14736	=>	65127,
		14737	=>	65127,
		14738	=>	65128,
		14739	=>	65128,
		14740	=>	65129,
		14741	=>	65129,
		14742	=>	65130,
		14743	=>	65130,
		14744	=>	65131,
		14745	=>	65131,
		14746	=>	65132,
		14747	=>	65132,
		14748	=>	65133,
		14749	=>	65133,
		14750	=>	65134,
		14751	=>	65134,
		14752	=>	65135,
		14753	=>	65135,
		14754	=>	65136,
		14755	=>	65136,
		14756	=>	65137,
		14757	=>	65137,
		14758	=>	65138,
		14759	=>	65138,
		14760	=>	65139,
		14761	=>	65139,
		14762	=>	65140,
		14763	=>	65140,
		14764	=>	65141,
		14765	=>	65141,
		14766	=>	65142,
		14767	=>	65142,
		14768	=>	65143,
		14769	=>	65143,
		14770	=>	65143,
		14771	=>	65144,
		14772	=>	65144,
		14773	=>	65145,
		14774	=>	65145,
		14775	=>	65146,
		14776	=>	65146,
		14777	=>	65147,
		14778	=>	65147,
		14779	=>	65148,
		14780	=>	65148,
		14781	=>	65149,
		14782	=>	65149,
		14783	=>	65150,
		14784	=>	65150,
		14785	=>	65151,
		14786	=>	65151,
		14787	=>	65152,
		14788	=>	65152,
		14789	=>	65153,
		14790	=>	65153,
		14791	=>	65154,
		14792	=>	65154,
		14793	=>	65155,
		14794	=>	65155,
		14795	=>	65155,
		14796	=>	65156,
		14797	=>	65156,
		14798	=>	65157,
		14799	=>	65157,
		14800	=>	65158,
		14801	=>	65158,
		14802	=>	65159,
		14803	=>	65159,
		14804	=>	65160,
		14805	=>	65160,
		14806	=>	65161,
		14807	=>	65161,
		14808	=>	65162,
		14809	=>	65162,
		14810	=>	65163,
		14811	=>	65163,
		14812	=>	65164,
		14813	=>	65164,
		14814	=>	65164,
		14815	=>	65165,
		14816	=>	65165,
		14817	=>	65166,
		14818	=>	65166,
		14819	=>	65167,
		14820	=>	65167,
		14821	=>	65168,
		14822	=>	65168,
		14823	=>	65169,
		14824	=>	65169,
		14825	=>	65170,
		14826	=>	65170,
		14827	=>	65171,
		14828	=>	65171,
		14829	=>	65172,
		14830	=>	65172,
		14831	=>	65172,
		14832	=>	65173,
		14833	=>	65173,
		14834	=>	65174,
		14835	=>	65174,
		14836	=>	65175,
		14837	=>	65175,
		14838	=>	65176,
		14839	=>	65176,
		14840	=>	65177,
		14841	=>	65177,
		14842	=>	65178,
		14843	=>	65178,
		14844	=>	65178,
		14845	=>	65179,
		14846	=>	65179,
		14847	=>	65180,
		14848	=>	65180,
		14849	=>	65181,
		14850	=>	65181,
		14851	=>	65182,
		14852	=>	65182,
		14853	=>	65183,
		14854	=>	65183,
		14855	=>	65184,
		14856	=>	65184,
		14857	=>	65184,
		14858	=>	65185,
		14859	=>	65185,
		14860	=>	65186,
		14861	=>	65186,
		14862	=>	65187,
		14863	=>	65187,
		14864	=>	65188,
		14865	=>	65188,
		14866	=>	65189,
		14867	=>	65189,
		14868	=>	65190,
		14869	=>	65190,
		14870	=>	65190,
		14871	=>	65191,
		14872	=>	65191,
		14873	=>	65192,
		14874	=>	65192,
		14875	=>	65193,
		14876	=>	65193,
		14877	=>	65194,
		14878	=>	65194,
		14879	=>	65194,
		14880	=>	65195,
		14881	=>	65195,
		14882	=>	65196,
		14883	=>	65196,
		14884	=>	65197,
		14885	=>	65197,
		14886	=>	65198,
		14887	=>	65198,
		14888	=>	65199,
		14889	=>	65199,
		14890	=>	65199,
		14891	=>	65200,
		14892	=>	65200,
		14893	=>	65201,
		14894	=>	65201,
		14895	=>	65202,
		14896	=>	65202,
		14897	=>	65203,
		14898	=>	65203,
		14899	=>	65203,
		14900	=>	65204,
		14901	=>	65204,
		14902	=>	65205,
		14903	=>	65205,
		14904	=>	65206,
		14905	=>	65206,
		14906	=>	65207,
		14907	=>	65207,
		14908	=>	65207,
		14909	=>	65208,
		14910	=>	65208,
		14911	=>	65209,
		14912	=>	65209,
		14913	=>	65210,
		14914	=>	65210,
		14915	=>	65211,
		14916	=>	65211,
		14917	=>	65211,
		14918	=>	65212,
		14919	=>	65212,
		14920	=>	65213,
		14921	=>	65213,
		14922	=>	65214,
		14923	=>	65214,
		14924	=>	65215,
		14925	=>	65215,
		14926	=>	65215,
		14927	=>	65216,
		14928	=>	65216,
		14929	=>	65217,
		14930	=>	65217,
		14931	=>	65218,
		14932	=>	65218,
		14933	=>	65218,
		14934	=>	65219,
		14935	=>	65219,
		14936	=>	65220,
		14937	=>	65220,
		14938	=>	65221,
		14939	=>	65221,
		14940	=>	65221,
		14941	=>	65222,
		14942	=>	65222,
		14943	=>	65223,
		14944	=>	65223,
		14945	=>	65224,
		14946	=>	65224,
		14947	=>	65225,
		14948	=>	65225,
		14949	=>	65225,
		14950	=>	65226,
		14951	=>	65226,
		14952	=>	65227,
		14953	=>	65227,
		14954	=>	65228,
		14955	=>	65228,
		14956	=>	65228,
		14957	=>	65229,
		14958	=>	65229,
		14959	=>	65230,
		14960	=>	65230,
		14961	=>	65231,
		14962	=>	65231,
		14963	=>	65231,
		14964	=>	65232,
		14965	=>	65232,
		14966	=>	65233,
		14967	=>	65233,
		14968	=>	65234,
		14969	=>	65234,
		14970	=>	65234,
		14971	=>	65235,
		14972	=>	65235,
		14973	=>	65236,
		14974	=>	65236,
		14975	=>	65236,
		14976	=>	65237,
		14977	=>	65237,
		14978	=>	65238,
		14979	=>	65238,
		14980	=>	65239,
		14981	=>	65239,
		14982	=>	65239,
		14983	=>	65240,
		14984	=>	65240,
		14985	=>	65241,
		14986	=>	65241,
		14987	=>	65242,
		14988	=>	65242,
		14989	=>	65242,
		14990	=>	65243,
		14991	=>	65243,
		14992	=>	65244,
		14993	=>	65244,
		14994	=>	65244,
		14995	=>	65245,
		14996	=>	65245,
		14997	=>	65246,
		14998	=>	65246,
		14999	=>	65247,
		15000	=>	65247,
		15001	=>	65247,
		15002	=>	65248,
		15003	=>	65248,
		15004	=>	65249,
		15005	=>	65249,
		15006	=>	65249,
		15007	=>	65250,
		15008	=>	65250,
		15009	=>	65251,
		15010	=>	65251,
		15011	=>	65252,
		15012	=>	65252,
		15013	=>	65252,
		15014	=>	65253,
		15015	=>	65253,
		15016	=>	65254,
		15017	=>	65254,
		15018	=>	65254,
		15019	=>	65255,
		15020	=>	65255,
		15021	=>	65256,
		15022	=>	65256,
		15023	=>	65256,
		15024	=>	65257,
		15025	=>	65257,
		15026	=>	65258,
		15027	=>	65258,
		15028	=>	65258,
		15029	=>	65259,
		15030	=>	65259,
		15031	=>	65260,
		15032	=>	65260,
		15033	=>	65261,
		15034	=>	65261,
		15035	=>	65261,
		15036	=>	65262,
		15037	=>	65262,
		15038	=>	65263,
		15039	=>	65263,
		15040	=>	65263,
		15041	=>	65264,
		15042	=>	65264,
		15043	=>	65265,
		15044	=>	65265,
		15045	=>	65265,
		15046	=>	65266,
		15047	=>	65266,
		15048	=>	65267,
		15049	=>	65267,
		15050	=>	65267,
		15051	=>	65268,
		15052	=>	65268,
		15053	=>	65269,
		15054	=>	65269,
		15055	=>	65269,
		15056	=>	65270,
		15057	=>	65270,
		15058	=>	65271,
		15059	=>	65271,
		15060	=>	65271,
		15061	=>	65272,
		15062	=>	65272,
		15063	=>	65273,
		15064	=>	65273,
		15065	=>	65273,
		15066	=>	65274,
		15067	=>	65274,
		15068	=>	65275,
		15069	=>	65275,
		15070	=>	65275,
		15071	=>	65276,
		15072	=>	65276,
		15073	=>	65277,
		15074	=>	65277,
		15075	=>	65277,
		15076	=>	65278,
		15077	=>	65278,
		15078	=>	65278,
		15079	=>	65279,
		15080	=>	65279,
		15081	=>	65280,
		15082	=>	65280,
		15083	=>	65280,
		15084	=>	65281,
		15085	=>	65281,
		15086	=>	65282,
		15087	=>	65282,
		15088	=>	65282,
		15089	=>	65283,
		15090	=>	65283,
		15091	=>	65284,
		15092	=>	65284,
		15093	=>	65284,
		15094	=>	65285,
		15095	=>	65285,
		15096	=>	65285,
		15097	=>	65286,
		15098	=>	65286,
		15099	=>	65287,
		15100	=>	65287,
		15101	=>	65287,
		15102	=>	65288,
		15103	=>	65288,
		15104	=>	65289,
		15105	=>	65289,
		15106	=>	65289,
		15107	=>	65290,
		15108	=>	65290,
		15109	=>	65290,
		15110	=>	65291,
		15111	=>	65291,
		15112	=>	65292,
		15113	=>	65292,
		15114	=>	65292,
		15115	=>	65293,
		15116	=>	65293,
		15117	=>	65294,
		15118	=>	65294,
		15119	=>	65294,
		15120	=>	65295,
		15121	=>	65295,
		15122	=>	65295,
		15123	=>	65296,
		15124	=>	65296,
		15125	=>	65297,
		15126	=>	65297,
		15127	=>	65297,
		15128	=>	65298,
		15129	=>	65298,
		15130	=>	65298,
		15131	=>	65299,
		15132	=>	65299,
		15133	=>	65300,
		15134	=>	65300,
		15135	=>	65300,
		15136	=>	65301,
		15137	=>	65301,
		15138	=>	65301,
		15139	=>	65302,
		15140	=>	65302,
		15141	=>	65303,
		15142	=>	65303,
		15143	=>	65303,
		15144	=>	65304,
		15145	=>	65304,
		15146	=>	65304,
		15147	=>	65305,
		15148	=>	65305,
		15149	=>	65306,
		15150	=>	65306,
		15151	=>	65306,
		15152	=>	65307,
		15153	=>	65307,
		15154	=>	65307,
		15155	=>	65308,
		15156	=>	65308,
		15157	=>	65309,
		15158	=>	65309,
		15159	=>	65309,
		15160	=>	65310,
		15161	=>	65310,
		15162	=>	65310,
		15163	=>	65311,
		15164	=>	65311,
		15165	=>	65311,
		15166	=>	65312,
		15167	=>	65312,
		15168	=>	65313,
		15169	=>	65313,
		15170	=>	65313,
		15171	=>	65314,
		15172	=>	65314,
		15173	=>	65314,
		15174	=>	65315,
		15175	=>	65315,
		15176	=>	65315,
		15177	=>	65316,
		15178	=>	65316,
		15179	=>	65317,
		15180	=>	65317,
		15181	=>	65317,
		15182	=>	65318,
		15183	=>	65318,
		15184	=>	65318,
		15185	=>	65319,
		15186	=>	65319,
		15187	=>	65319,
		15188	=>	65320,
		15189	=>	65320,
		15190	=>	65321,
		15191	=>	65321,
		15192	=>	65321,
		15193	=>	65322,
		15194	=>	65322,
		15195	=>	65322,
		15196	=>	65323,
		15197	=>	65323,
		15198	=>	65323,
		15199	=>	65324,
		15200	=>	65324,
		15201	=>	65324,
		15202	=>	65325,
		15203	=>	65325,
		15204	=>	65326,
		15205	=>	65326,
		15206	=>	65326,
		15207	=>	65327,
		15208	=>	65327,
		15209	=>	65327,
		15210	=>	65328,
		15211	=>	65328,
		15212	=>	65328,
		15213	=>	65329,
		15214	=>	65329,
		15215	=>	65329,
		15216	=>	65330,
		15217	=>	65330,
		15218	=>	65330,
		15219	=>	65331,
		15220	=>	65331,
		15221	=>	65332,
		15222	=>	65332,
		15223	=>	65332,
		15224	=>	65333,
		15225	=>	65333,
		15226	=>	65333,
		15227	=>	65334,
		15228	=>	65334,
		15229	=>	65334,
		15230	=>	65335,
		15231	=>	65335,
		15232	=>	65335,
		15233	=>	65336,
		15234	=>	65336,
		15235	=>	65336,
		15236	=>	65337,
		15237	=>	65337,
		15238	=>	65337,
		15239	=>	65338,
		15240	=>	65338,
		15241	=>	65338,
		15242	=>	65339,
		15243	=>	65339,
		15244	=>	65339,
		15245	=>	65340,
		15246	=>	65340,
		15247	=>	65341,
		15248	=>	65341,
		15249	=>	65341,
		15250	=>	65342,
		15251	=>	65342,
		15252	=>	65342,
		15253	=>	65343,
		15254	=>	65343,
		15255	=>	65343,
		15256	=>	65344,
		15257	=>	65344,
		15258	=>	65344,
		15259	=>	65345,
		15260	=>	65345,
		15261	=>	65345,
		15262	=>	65346,
		15263	=>	65346,
		15264	=>	65346,
		15265	=>	65347,
		15266	=>	65347,
		15267	=>	65347,
		15268	=>	65348,
		15269	=>	65348,
		15270	=>	65348,
		15271	=>	65349,
		15272	=>	65349,
		15273	=>	65349,
		15274	=>	65350,
		15275	=>	65350,
		15276	=>	65350,
		15277	=>	65351,
		15278	=>	65351,
		15279	=>	65351,
		15280	=>	65352,
		15281	=>	65352,
		15282	=>	65352,
		15283	=>	65353,
		15284	=>	65353,
		15285	=>	65353,
		15286	=>	65354,
		15287	=>	65354,
		15288	=>	65354,
		15289	=>	65355,
		15290	=>	65355,
		15291	=>	65355,
		15292	=>	65356,
		15293	=>	65356,
		15294	=>	65356,
		15295	=>	65357,
		15296	=>	65357,
		15297	=>	65357,
		15298	=>	65358,
		15299	=>	65358,
		15300	=>	65358,
		15301	=>	65359,
		15302	=>	65359,
		15303	=>	65359,
		15304	=>	65360,
		15305	=>	65360,
		15306	=>	65360,
		15307	=>	65360,
		15308	=>	65361,
		15309	=>	65361,
		15310	=>	65361,
		15311	=>	65362,
		15312	=>	65362,
		15313	=>	65362,
		15314	=>	65363,
		15315	=>	65363,
		15316	=>	65363,
		15317	=>	65364,
		15318	=>	65364,
		15319	=>	65364,
		15320	=>	65365,
		15321	=>	65365,
		15322	=>	65365,
		15323	=>	65366,
		15324	=>	65366,
		15325	=>	65366,
		15326	=>	65367,
		15327	=>	65367,
		15328	=>	65367,
		15329	=>	65368,
		15330	=>	65368,
		15331	=>	65368,
		15332	=>	65368,
		15333	=>	65369,
		15334	=>	65369,
		15335	=>	65369,
		15336	=>	65370,
		15337	=>	65370,
		15338	=>	65370,
		15339	=>	65371,
		15340	=>	65371,
		15341	=>	65371,
		15342	=>	65372,
		15343	=>	65372,
		15344	=>	65372,
		15345	=>	65373,
		15346	=>	65373,
		15347	=>	65373,
		15348	=>	65373,
		15349	=>	65374,
		15350	=>	65374,
		15351	=>	65374,
		15352	=>	65375,
		15353	=>	65375,
		15354	=>	65375,
		15355	=>	65376,
		15356	=>	65376,
		15357	=>	65376,
		15358	=>	65377,
		15359	=>	65377,
		15360	=>	65377,
		15361	=>	65378,
		15362	=>	65378,
		15363	=>	65378,
		15364	=>	65378,
		15365	=>	65379,
		15366	=>	65379,
		15367	=>	65379,
		15368	=>	65380,
		15369	=>	65380,
		15370	=>	65380,
		15371	=>	65381,
		15372	=>	65381,
		15373	=>	65381,
		15374	=>	65381,
		15375	=>	65382,
		15376	=>	65382,
		15377	=>	65382,
		15378	=>	65383,
		15379	=>	65383,
		15380	=>	65383,
		15381	=>	65384,
		15382	=>	65384,
		15383	=>	65384,
		15384	=>	65385,
		15385	=>	65385,
		15386	=>	65385,
		15387	=>	65385,
		15388	=>	65386,
		15389	=>	65386,
		15390	=>	65386,
		15391	=>	65387,
		15392	=>	65387,
		15393	=>	65387,
		15394	=>	65388,
		15395	=>	65388,
		15396	=>	65388,
		15397	=>	65388,
		15398	=>	65389,
		15399	=>	65389,
		15400	=>	65389,
		15401	=>	65390,
		15402	=>	65390,
		15403	=>	65390,
		15404	=>	65390,
		15405	=>	65391,
		15406	=>	65391,
		15407	=>	65391,
		15408	=>	65392,
		15409	=>	65392,
		15410	=>	65392,
		15411	=>	65393,
		15412	=>	65393,
		15413	=>	65393,
		15414	=>	65393,
		15415	=>	65394,
		15416	=>	65394,
		15417	=>	65394,
		15418	=>	65395,
		15419	=>	65395,
		15420	=>	65395,
		15421	=>	65395,
		15422	=>	65396,
		15423	=>	65396,
		15424	=>	65396,
		15425	=>	65397,
		15426	=>	65397,
		15427	=>	65397,
		15428	=>	65397,
		15429	=>	65398,
		15430	=>	65398,
		15431	=>	65398,
		15432	=>	65399,
		15433	=>	65399,
		15434	=>	65399,
		15435	=>	65399,
		15436	=>	65400,
		15437	=>	65400,
		15438	=>	65400,
		15439	=>	65401,
		15440	=>	65401,
		15441	=>	65401,
		15442	=>	65401,
		15443	=>	65402,
		15444	=>	65402,
		15445	=>	65402,
		15446	=>	65403,
		15447	=>	65403,
		15448	=>	65403,
		15449	=>	65403,
		15450	=>	65404,
		15451	=>	65404,
		15452	=>	65404,
		15453	=>	65405,
		15454	=>	65405,
		15455	=>	65405,
		15456	=>	65405,
		15457	=>	65406,
		15458	=>	65406,
		15459	=>	65406,
		15460	=>	65407,
		15461	=>	65407,
		15462	=>	65407,
		15463	=>	65407,
		15464	=>	65408,
		15465	=>	65408,
		15466	=>	65408,
		15467	=>	65408,
		15468	=>	65409,
		15469	=>	65409,
		15470	=>	65409,
		15471	=>	65410,
		15472	=>	65410,
		15473	=>	65410,
		15474	=>	65410,
		15475	=>	65411,
		15476	=>	65411,
		15477	=>	65411,
		15478	=>	65411,
		15479	=>	65412,
		15480	=>	65412,
		15481	=>	65412,
		15482	=>	65413,
		15483	=>	65413,
		15484	=>	65413,
		15485	=>	65413,
		15486	=>	65414,
		15487	=>	65414,
		15488	=>	65414,
		15489	=>	65414,
		15490	=>	65415,
		15491	=>	65415,
		15492	=>	65415,
		15493	=>	65416,
		15494	=>	65416,
		15495	=>	65416,
		15496	=>	65416,
		15497	=>	65417,
		15498	=>	65417,
		15499	=>	65417,
		15500	=>	65417,
		15501	=>	65418,
		15502	=>	65418,
		15503	=>	65418,
		15504	=>	65418,
		15505	=>	65419,
		15506	=>	65419,
		15507	=>	65419,
		15508	=>	65420,
		15509	=>	65420,
		15510	=>	65420,
		15511	=>	65420,
		15512	=>	65421,
		15513	=>	65421,
		15514	=>	65421,
		15515	=>	65421,
		15516	=>	65422,
		15517	=>	65422,
		15518	=>	65422,
		15519	=>	65422,
		15520	=>	65423,
		15521	=>	65423,
		15522	=>	65423,
		15523	=>	65423,
		15524	=>	65424,
		15525	=>	65424,
		15526	=>	65424,
		15527	=>	65424,
		15528	=>	65425,
		15529	=>	65425,
		15530	=>	65425,
		15531	=>	65425,
		15532	=>	65426,
		15533	=>	65426,
		15534	=>	65426,
		15535	=>	65427,
		15536	=>	65427,
		15537	=>	65427,
		15538	=>	65427,
		15539	=>	65428,
		15540	=>	65428,
		15541	=>	65428,
		15542	=>	65428,
		15543	=>	65429,
		15544	=>	65429,
		15545	=>	65429,
		15546	=>	65429,
		15547	=>	65430,
		15548	=>	65430,
		15549	=>	65430,
		15550	=>	65430,
		15551	=>	65431,
		15552	=>	65431,
		15553	=>	65431,
		15554	=>	65431,
		15555	=>	65432,
		15556	=>	65432,
		15557	=>	65432,
		15558	=>	65432,
		15559	=>	65433,
		15560	=>	65433,
		15561	=>	65433,
		15562	=>	65433,
		15563	=>	65434,
		15564	=>	65434,
		15565	=>	65434,
		15566	=>	65434,
		15567	=>	65435,
		15568	=>	65435,
		15569	=>	65435,
		15570	=>	65435,
		15571	=>	65436,
		15572	=>	65436,
		15573	=>	65436,
		15574	=>	65436,
		15575	=>	65436,
		15576	=>	65437,
		15577	=>	65437,
		15578	=>	65437,
		15579	=>	65437,
		15580	=>	65438,
		15581	=>	65438,
		15582	=>	65438,
		15583	=>	65438,
		15584	=>	65439,
		15585	=>	65439,
		15586	=>	65439,
		15587	=>	65439,
		15588	=>	65440,
		15589	=>	65440,
		15590	=>	65440,
		15591	=>	65440,
		15592	=>	65441,
		15593	=>	65441,
		15594	=>	65441,
		15595	=>	65441,
		15596	=>	65442,
		15597	=>	65442,
		15598	=>	65442,
		15599	=>	65442,
		15600	=>	65442,
		15601	=>	65443,
		15602	=>	65443,
		15603	=>	65443,
		15604	=>	65443,
		15605	=>	65444,
		15606	=>	65444,
		15607	=>	65444,
		15608	=>	65444,
		15609	=>	65445,
		15610	=>	65445,
		15611	=>	65445,
		15612	=>	65445,
		15613	=>	65446,
		15614	=>	65446,
		15615	=>	65446,
		15616	=>	65446,
		15617	=>	65446,
		15618	=>	65447,
		15619	=>	65447,
		15620	=>	65447,
		15621	=>	65447,
		15622	=>	65448,
		15623	=>	65448,
		15624	=>	65448,
		15625	=>	65448,
		15626	=>	65449,
		15627	=>	65449,
		15628	=>	65449,
		15629	=>	65449,
		15630	=>	65449,
		15631	=>	65450,
		15632	=>	65450,
		15633	=>	65450,
		15634	=>	65450,
		15635	=>	65451,
		15636	=>	65451,
		15637	=>	65451,
		15638	=>	65451,
		15639	=>	65451,
		15640	=>	65452,
		15641	=>	65452,
		15642	=>	65452,
		15643	=>	65452,
		15644	=>	65453,
		15645	=>	65453,
		15646	=>	65453,
		15647	=>	65453,
		15648	=>	65453,
		15649	=>	65454,
		15650	=>	65454,
		15651	=>	65454,
		15652	=>	65454,
		15653	=>	65455,
		15654	=>	65455,
		15655	=>	65455,
		15656	=>	65455,
		15657	=>	65455,
		15658	=>	65456,
		15659	=>	65456,
		15660	=>	65456,
		15661	=>	65456,
		15662	=>	65457,
		15663	=>	65457,
		15664	=>	65457,
		15665	=>	65457,
		15666	=>	65457,
		15667	=>	65458,
		15668	=>	65458,
		15669	=>	65458,
		15670	=>	65458,
		15671	=>	65458,
		15672	=>	65459,
		15673	=>	65459,
		15674	=>	65459,
		15675	=>	65459,
		15676	=>	65460,
		15677	=>	65460,
		15678	=>	65460,
		15679	=>	65460,
		15680	=>	65460,
		15681	=>	65461,
		15682	=>	65461,
		15683	=>	65461,
		15684	=>	65461,
		15685	=>	65461,
		15686	=>	65462,
		15687	=>	65462,
		15688	=>	65462,
		15689	=>	65462,
		15690	=>	65462,
		15691	=>	65463,
		15692	=>	65463,
		15693	=>	65463,
		15694	=>	65463,
		15695	=>	65464,
		15696	=>	65464,
		15697	=>	65464,
		15698	=>	65464,
		15699	=>	65464,
		15700	=>	65465,
		15701	=>	65465,
		15702	=>	65465,
		15703	=>	65465,
		15704	=>	65465,
		15705	=>	65466,
		15706	=>	65466,
		15707	=>	65466,
		15708	=>	65466,
		15709	=>	65466,
		15710	=>	65467,
		15711	=>	65467,
		15712	=>	65467,
		15713	=>	65467,
		15714	=>	65467,
		15715	=>	65468,
		15716	=>	65468,
		15717	=>	65468,
		15718	=>	65468,
		15719	=>	65468,
		15720	=>	65469,
		15721	=>	65469,
		15722	=>	65469,
		15723	=>	65469,
		15724	=>	65469,
		15725	=>	65470,
		15726	=>	65470,
		15727	=>	65470,
		15728	=>	65470,
		15729	=>	65470,
		15730	=>	65471,
		15731	=>	65471,
		15732	=>	65471,
		15733	=>	65471,
		15734	=>	65471,
		15735	=>	65472,
		15736	=>	65472,
		15737	=>	65472,
		15738	=>	65472,
		15739	=>	65472,
		15740	=>	65473,
		15741	=>	65473,
		15742	=>	65473,
		15743	=>	65473,
		15744	=>	65473,
		15745	=>	65474,
		15746	=>	65474,
		15747	=>	65474,
		15748	=>	65474,
		15749	=>	65474,
		15750	=>	65474,
		15751	=>	65475,
		15752	=>	65475,
		15753	=>	65475,
		15754	=>	65475,
		15755	=>	65475,
		15756	=>	65476,
		15757	=>	65476,
		15758	=>	65476,
		15759	=>	65476,
		15760	=>	65476,
		15761	=>	65477,
		15762	=>	65477,
		15763	=>	65477,
		15764	=>	65477,
		15765	=>	65477,
		15766	=>	65478,
		15767	=>	65478,
		15768	=>	65478,
		15769	=>	65478,
		15770	=>	65478,
		15771	=>	65478,
		15772	=>	65479,
		15773	=>	65479,
		15774	=>	65479,
		15775	=>	65479,
		15776	=>	65479,
		15777	=>	65480,
		15778	=>	65480,
		15779	=>	65480,
		15780	=>	65480,
		15781	=>	65480,
		15782	=>	65480,
		15783	=>	65481,
		15784	=>	65481,
		15785	=>	65481,
		15786	=>	65481,
		15787	=>	65481,
		15788	=>	65482,
		15789	=>	65482,
		15790	=>	65482,
		15791	=>	65482,
		15792	=>	65482,
		15793	=>	65482,
		15794	=>	65483,
		15795	=>	65483,
		15796	=>	65483,
		15797	=>	65483,
		15798	=>	65483,
		15799	=>	65483,
		15800	=>	65484,
		15801	=>	65484,
		15802	=>	65484,
		15803	=>	65484,
		15804	=>	65484,
		15805	=>	65485,
		15806	=>	65485,
		15807	=>	65485,
		15808	=>	65485,
		15809	=>	65485,
		15810	=>	65485,
		15811	=>	65486,
		15812	=>	65486,
		15813	=>	65486,
		15814	=>	65486,
		15815	=>	65486,
		15816	=>	65486,
		15817	=>	65487,
		15818	=>	65487,
		15819	=>	65487,
		15820	=>	65487,
		15821	=>	65487,
		15822	=>	65487,
		15823	=>	65488,
		15824	=>	65488,
		15825	=>	65488,
		15826	=>	65488,
		15827	=>	65488,
		15828	=>	65488,
		15829	=>	65489,
		15830	=>	65489,
		15831	=>	65489,
		15832	=>	65489,
		15833	=>	65489,
		15834	=>	65489,
		15835	=>	65490,
		15836	=>	65490,
		15837	=>	65490,
		15838	=>	65490,
		15839	=>	65490,
		15840	=>	65490,
		15841	=>	65491,
		15842	=>	65491,
		15843	=>	65491,
		15844	=>	65491,
		15845	=>	65491,
		15846	=>	65491,
		15847	=>	65492,
		15848	=>	65492,
		15849	=>	65492,
		15850	=>	65492,
		15851	=>	65492,
		15852	=>	65492,
		15853	=>	65493,
		15854	=>	65493,
		15855	=>	65493,
		15856	=>	65493,
		15857	=>	65493,
		15858	=>	65493,
		15859	=>	65494,
		15860	=>	65494,
		15861	=>	65494,
		15862	=>	65494,
		15863	=>	65494,
		15864	=>	65494,
		15865	=>	65494,
		15866	=>	65495,
		15867	=>	65495,
		15868	=>	65495,
		15869	=>	65495,
		15870	=>	65495,
		15871	=>	65495,
		15872	=>	65496,
		15873	=>	65496,
		15874	=>	65496,
		15875	=>	65496,
		15876	=>	65496,
		15877	=>	65496,
		15878	=>	65496,
		15879	=>	65497,
		15880	=>	65497,
		15881	=>	65497,
		15882	=>	65497,
		15883	=>	65497,
		15884	=>	65497,
		15885	=>	65498,
		15886	=>	65498,
		15887	=>	65498,
		15888	=>	65498,
		15889	=>	65498,
		15890	=>	65498,
		15891	=>	65498,
		15892	=>	65499,
		15893	=>	65499,
		15894	=>	65499,
		15895	=>	65499,
		15896	=>	65499,
		15897	=>	65499,
		15898	=>	65499,
		15899	=>	65500,
		15900	=>	65500,
		15901	=>	65500,
		15902	=>	65500,
		15903	=>	65500,
		15904	=>	65500,
		15905	=>	65500,
		15906	=>	65501,
		15907	=>	65501,
		15908	=>	65501,
		15909	=>	65501,
		15910	=>	65501,
		15911	=>	65501,
		15912	=>	65501,
		15913	=>	65502,
		15914	=>	65502,
		15915	=>	65502,
		15916	=>	65502,
		15917	=>	65502,
		15918	=>	65502,
		15919	=>	65502,
		15920	=>	65503,
		15921	=>	65503,
		15922	=>	65503,
		15923	=>	65503,
		15924	=>	65503,
		15925	=>	65503,
		15926	=>	65503,
		15927	=>	65504,
		15928	=>	65504,
		15929	=>	65504,
		15930	=>	65504,
		15931	=>	65504,
		15932	=>	65504,
		15933	=>	65504,
		15934	=>	65505,
		15935	=>	65505,
		15936	=>	65505,
		15937	=>	65505,
		15938	=>	65505,
		15939	=>	65505,
		15940	=>	65505,
		15941	=>	65505,
		15942	=>	65506,
		15943	=>	65506,
		15944	=>	65506,
		15945	=>	65506,
		15946	=>	65506,
		15947	=>	65506,
		15948	=>	65506,
		15949	=>	65507,
		15950	=>	65507,
		15951	=>	65507,
		15952	=>	65507,
		15953	=>	65507,
		15954	=>	65507,
		15955	=>	65507,
		15956	=>	65507,
		15957	=>	65508,
		15958	=>	65508,
		15959	=>	65508,
		15960	=>	65508,
		15961	=>	65508,
		15962	=>	65508,
		15963	=>	65508,
		15964	=>	65508,
		15965	=>	65509,
		15966	=>	65509,
		15967	=>	65509,
		15968	=>	65509,
		15969	=>	65509,
		15970	=>	65509,
		15971	=>	65509,
		15972	=>	65509,
		15973	=>	65510,
		15974	=>	65510,
		15975	=>	65510,
		15976	=>	65510,
		15977	=>	65510,
		15978	=>	65510,
		15979	=>	65510,
		15980	=>	65510,
		15981	=>	65511,
		15982	=>	65511,
		15983	=>	65511,
		15984	=>	65511,
		15985	=>	65511,
		15986	=>	65511,
		15987	=>	65511,
		15988	=>	65511,
		15989	=>	65512,
		15990	=>	65512,
		15991	=>	65512,
		15992	=>	65512,
		15993	=>	65512,
		15994	=>	65512,
		15995	=>	65512,
		15996	=>	65512,
		15997	=>	65512,
		15998	=>	65513,
		15999	=>	65513,
		16000	=>	65513,
		16001	=>	65513,
		16002	=>	65513,
		16003	=>	65513,
		16004	=>	65513,
		16005	=>	65513,
		16006	=>	65513,
		16007	=>	65514,
		16008	=>	65514,
		16009	=>	65514,
		16010	=>	65514,
		16011	=>	65514,
		16012	=>	65514,
		16013	=>	65514,
		16014	=>	65514,
		16015	=>	65514,
		16016	=>	65515,
		16017	=>	65515,
		16018	=>	65515,
		16019	=>	65515,
		16020	=>	65515,
		16021	=>	65515,
		16022	=>	65515,
		16023	=>	65515,
		16024	=>	65515,
		16025	=>	65516,
		16026	=>	65516,
		16027	=>	65516,
		16028	=>	65516,
		16029	=>	65516,
		16030	=>	65516,
		16031	=>	65516,
		16032	=>	65516,
		16033	=>	65516,
		16034	=>	65517,
		16035	=>	65517,
		16036	=>	65517,
		16037	=>	65517,
		16038	=>	65517,
		16039	=>	65517,
		16040	=>	65517,
		16041	=>	65517,
		16042	=>	65517,
		16043	=>	65517,
		16044	=>	65518,
		16045	=>	65518,
		16046	=>	65518,
		16047	=>	65518,
		16048	=>	65518,
		16049	=>	65518,
		16050	=>	65518,
		16051	=>	65518,
		16052	=>	65518,
		16053	=>	65519,
		16054	=>	65519,
		16055	=>	65519,
		16056	=>	65519,
		16057	=>	65519,
		16058	=>	65519,
		16059	=>	65519,
		16060	=>	65519,
		16061	=>	65519,
		16062	=>	65519,
		16063	=>	65519,
		16064	=>	65520,
		16065	=>	65520,
		16066	=>	65520,
		16067	=>	65520,
		16068	=>	65520,
		16069	=>	65520,
		16070	=>	65520,
		16071	=>	65520,
		16072	=>	65520,
		16073	=>	65520,
		16074	=>	65521,
		16075	=>	65521,
		16076	=>	65521,
		16077	=>	65521,
		16078	=>	65521,
		16079	=>	65521,
		16080	=>	65521,
		16081	=>	65521,
		16082	=>	65521,
		16083	=>	65521,
		16084	=>	65521,
		16085	=>	65522,
		16086	=>	65522,
		16087	=>	65522,
		16088	=>	65522,
		16089	=>	65522,
		16090	=>	65522,
		16091	=>	65522,
		16092	=>	65522,
		16093	=>	65522,
		16094	=>	65522,
		16095	=>	65522,
		16096	=>	65523,
		16097	=>	65523,
		16098	=>	65523,
		16099	=>	65523,
		16100	=>	65523,
		16101	=>	65523,
		16102	=>	65523,
		16103	=>	65523,
		16104	=>	65523,
		16105	=>	65523,
		16106	=>	65523,
		16107	=>	65523,
		16108	=>	65524,
		16109	=>	65524,
		16110	=>	65524,
		16111	=>	65524,
		16112	=>	65524,
		16113	=>	65524,
		16114	=>	65524,
		16115	=>	65524,
		16116	=>	65524,
		16117	=>	65524,
		16118	=>	65524,
		16119	=>	65524,
		16120	=>	65525,
		16121	=>	65525,
		16122	=>	65525,
		16123	=>	65525,
		16124	=>	65525,
		16125	=>	65525,
		16126	=>	65525,
		16127	=>	65525,
		16128	=>	65525,
		16129	=>	65525,
		16130	=>	65525,
		16131	=>	65525,
		16132	=>	65525,
		16133	=>	65526,
		16134	=>	65526,
		16135	=>	65526,
		16136	=>	65526,
		16137	=>	65526,
		16138	=>	65526,
		16139	=>	65526,
		16140	=>	65526,
		16141	=>	65526,
		16142	=>	65526,
		16143	=>	65526,
		16144	=>	65526,
		16145	=>	65526,
		16146	=>	65526,
		16147	=>	65527,
		16148	=>	65527,
		16149	=>	65527,
		16150	=>	65527,
		16151	=>	65527,
		16152	=>	65527,
		16153	=>	65527,
		16154	=>	65527,
		16155	=>	65527,
		16156	=>	65527,
		16157	=>	65527,
		16158	=>	65527,
		16159	=>	65527,
		16160	=>	65527,
		16161	=>	65528,
		16162	=>	65528,
		16163	=>	65528,
		16164	=>	65528,
		16165	=>	65528,
		16166	=>	65528,
		16167	=>	65528,
		16168	=>	65528,
		16169	=>	65528,
		16170	=>	65528,
		16171	=>	65528,
		16172	=>	65528,
		16173	=>	65528,
		16174	=>	65528,
		16175	=>	65528,
		16176	=>	65528,
		16177	=>	65529,
		16178	=>	65529,
		16179	=>	65529,
		16180	=>	65529,
		16181	=>	65529,
		16182	=>	65529,
		16183	=>	65529,
		16184	=>	65529,
		16185	=>	65529,
		16186	=>	65529,
		16187	=>	65529,
		16188	=>	65529,
		16189	=>	65529,
		16190	=>	65529,
		16191	=>	65529,
		16192	=>	65529,
		16193	=>	65530,
		16194	=>	65530,
		16195	=>	65530,
		16196	=>	65530,
		16197	=>	65530,
		16198	=>	65530,
		16199	=>	65530,
		16200	=>	65530,
		16201	=>	65530,
		16202	=>	65530,
		16203	=>	65530,
		16204	=>	65530,
		16205	=>	65530,
		16206	=>	65530,
		16207	=>	65530,
		16208	=>	65530,
		16209	=>	65530,
		16210	=>	65530,
		16211	=>	65530,
		16212	=>	65531,
		16213	=>	65531,
		16214	=>	65531,
		16215	=>	65531,
		16216	=>	65531,
		16217	=>	65531,
		16218	=>	65531,
		16219	=>	65531,
		16220	=>	65531,
		16221	=>	65531,
		16222	=>	65531,
		16223	=>	65531,
		16224	=>	65531,
		16225	=>	65531,
		16226	=>	65531,
		16227	=>	65531,
		16228	=>	65531,
		16229	=>	65531,
		16230	=>	65531,
		16231	=>	65531,
		16232	=>	65532,
		16233	=>	65532,
		16234	=>	65532,
		16235	=>	65532,
		16236	=>	65532,
		16237	=>	65532,
		16238	=>	65532,
		16239	=>	65532,
		16240	=>	65532,
		16241	=>	65532,
		16242	=>	65532,
		16243	=>	65532,
		16244	=>	65532,
		16245	=>	65532,
		16246	=>	65532,
		16247	=>	65532,
		16248	=>	65532,
		16249	=>	65532,
		16250	=>	65532,
		16251	=>	65532,
		16252	=>	65532,
		16253	=>	65532,
		16254	=>	65532,
		16255	=>	65532,
		16256	=>	65533,
		16257	=>	65533,
		16258	=>	65533,
		16259	=>	65533,
		16260	=>	65533,
		16261	=>	65533,
		16262	=>	65533,
		16263	=>	65533,
		16264	=>	65533,
		16265	=>	65533,
		16266	=>	65533,
		16267	=>	65533,
		16268	=>	65533,
		16269	=>	65533,
		16270	=>	65533,
		16271	=>	65533,
		16272	=>	65533,
		16273	=>	65533,
		16274	=>	65533,
		16275	=>	65533,
		16276	=>	65533,
		16277	=>	65533,
		16278	=>	65533,
		16279	=>	65533,
		16280	=>	65533,
		16281	=>	65533,
		16282	=>	65533,
		16283	=>	65533,
		16284	=>	65533,
		16285	=>	65534,
		16286	=>	65534,
		16287	=>	65534,
		16288	=>	65534,
		16289	=>	65534,
		16290	=>	65534,
		16291	=>	65534,
		16292	=>	65534,
		16293	=>	65534,
		16294	=>	65534,
		16295	=>	65534,
		16296	=>	65534,
		16297	=>	65534,
		16298	=>	65534,
		16299	=>	65534,
		16300	=>	65534,
		16301	=>	65534,
		16302	=>	65534,
		16303	=>	65534,
		16304	=>	65534,
		16305	=>	65534,
		16306	=>	65534,
		16307	=>	65534,
		16308	=>	65534,
		16309	=>	65534,
		16310	=>	65534,
		16311	=>	65534,
		16312	=>	65534,
		16313	=>	65534,
		16314	=>	65534,
		16315	=>	65534,
		16316	=>	65534,
		16317	=>	65534,
		16318	=>	65534,
		16319	=>	65534,
		16320	=>	65534,
		16321	=>	65534,
		16322	=>	65534,
		16323	=>	65534,
		16324	=>	65534,
		16325	=>	65534,
		16326	=>	65534,
		16327	=>	65535,
		16328	=>	65535,
		16329	=>	65535,
		16330	=>	65535,
		16331	=>	65535,
		16332	=>	65535,
		16333	=>	65535,
		16334	=>	65535,
		16335	=>	65535,
		16336	=>	65535,
		16337	=>	65535,
		16338	=>	65535,
		16339	=>	65535,
		16340	=>	65535,
		16341	=>	65535,
		16342	=>	65535,
		16343	=>	65535,
		16344	=>	65535,
		16345	=>	65535,
		16346	=>	65535,
		16347	=>	65535,
		16348	=>	65535,
		16349	=>	65535,
		16350	=>	65535,
		16351	=>	65535,
		16352	=>	65535,
		16353	=>	65535,
		16354	=>	65535,
		16355	=>	65535,
		16356	=>	65535,
		16357	=>	65535,
		16358	=>	65535,
		16359	=>	65535,
		16360	=>	65535,
		16361	=>	65535,
		16362	=>	65535,
		16363	=>	65535,
		16364	=>	65535,
		16365	=>	65535,
		16366	=>	65535,
		16367	=>	65535,
		16368	=>	65535,
		16369	=>	65535,
		16370	=>	65535,
		16371	=>	65535,
		16372	=>	65535,
		16373	=>	65535,
		16374	=>	65535,
		16375	=>	65535,
		16376	=>	65535,
		16377	=>	65535,
		16378	=>	65535,
		16379	=>	65535,
		16380	=>	65535,
		16381	=>	65535,
		16382	=>	65535,
		16383	=>	65535,
		16384	=>	65535,
		16385	=>	65535,
		16386	=>	65535,
		16387	=>	65535,
		16388	=>	65535,
		16389	=>	65535,
		16390	=>	65535,
		16391	=>	65535,
		16392	=>	65535,
		16393	=>	65535,
		16394	=>	65535,
		16395	=>	65535,
		16396	=>	65535,
		16397	=>	65535,
		16398	=>	65535,
		16399	=>	65535,
		16400	=>	65535,
		16401	=>	65535,
		16402	=>	65535,
		16403	=>	65535,
		16404	=>	65535,
		16405	=>	65535,
		16406	=>	65535,
		16407	=>	65535,
		16408	=>	65535,
		16409	=>	65535,
		16410	=>	65535,
		16411	=>	65535,
		16412	=>	65535,
		16413	=>	65535,
		16414	=>	65535,
		16415	=>	65535,
		16416	=>	65535,
		16417	=>	65535,
		16418	=>	65535,
		16419	=>	65535,
		16420	=>	65535,
		16421	=>	65535,
		16422	=>	65535,
		16423	=>	65535,
		16424	=>	65535,
		16425	=>	65535,
		16426	=>	65535,
		16427	=>	65535,
		16428	=>	65535,
		16429	=>	65535,
		16430	=>	65535,
		16431	=>	65535,
		16432	=>	65535,
		16433	=>	65535,
		16434	=>	65535,
		16435	=>	65535,
		16436	=>	65535,
		16437	=>	65535,
		16438	=>	65535,
		16439	=>	65535,
		16440	=>	65535,
		16441	=>	65535,
		16442	=>	65534,
		16443	=>	65534,
		16444	=>	65534,
		16445	=>	65534,
		16446	=>	65534,
		16447	=>	65534,
		16448	=>	65534,
		16449	=>	65534,
		16450	=>	65534,
		16451	=>	65534,
		16452	=>	65534,
		16453	=>	65534,
		16454	=>	65534,
		16455	=>	65534,
		16456	=>	65534,
		16457	=>	65534,
		16458	=>	65534,
		16459	=>	65534,
		16460	=>	65534,
		16461	=>	65534,
		16462	=>	65534,
		16463	=>	65534,
		16464	=>	65534,
		16465	=>	65534,
		16466	=>	65534,
		16467	=>	65534,
		16468	=>	65534,
		16469	=>	65534,
		16470	=>	65534,
		16471	=>	65534,
		16472	=>	65534,
		16473	=>	65534,
		16474	=>	65534,
		16475	=>	65534,
		16476	=>	65534,
		16477	=>	65534,
		16478	=>	65534,
		16479	=>	65534,
		16480	=>	65534,
		16481	=>	65534,
		16482	=>	65534,
		16483	=>	65534,
		16484	=>	65533,
		16485	=>	65533,
		16486	=>	65533,
		16487	=>	65533,
		16488	=>	65533,
		16489	=>	65533,
		16490	=>	65533,
		16491	=>	65533,
		16492	=>	65533,
		16493	=>	65533,
		16494	=>	65533,
		16495	=>	65533,
		16496	=>	65533,
		16497	=>	65533,
		16498	=>	65533,
		16499	=>	65533,
		16500	=>	65533,
		16501	=>	65533,
		16502	=>	65533,
		16503	=>	65533,
		16504	=>	65533,
		16505	=>	65533,
		16506	=>	65533,
		16507	=>	65533,
		16508	=>	65533,
		16509	=>	65533,
		16510	=>	65533,
		16511	=>	65533,
		16512	=>	65533,
		16513	=>	65532,
		16514	=>	65532,
		16515	=>	65532,
		16516	=>	65532,
		16517	=>	65532,
		16518	=>	65532,
		16519	=>	65532,
		16520	=>	65532,
		16521	=>	65532,
		16522	=>	65532,
		16523	=>	65532,
		16524	=>	65532,
		16525	=>	65532,
		16526	=>	65532,
		16527	=>	65532,
		16528	=>	65532,
		16529	=>	65532,
		16530	=>	65532,
		16531	=>	65532,
		16532	=>	65532,
		16533	=>	65532,
		16534	=>	65532,
		16535	=>	65532,
		16536	=>	65532,
		16537	=>	65531,
		16538	=>	65531,
		16539	=>	65531,
		16540	=>	65531,
		16541	=>	65531,
		16542	=>	65531,
		16543	=>	65531,
		16544	=>	65531,
		16545	=>	65531,
		16546	=>	65531,
		16547	=>	65531,
		16548	=>	65531,
		16549	=>	65531,
		16550	=>	65531,
		16551	=>	65531,
		16552	=>	65531,
		16553	=>	65531,
		16554	=>	65531,
		16555	=>	65531,
		16556	=>	65531,
		16557	=>	65530,
		16558	=>	65530,
		16559	=>	65530,
		16560	=>	65530,
		16561	=>	65530,
		16562	=>	65530,
		16563	=>	65530,
		16564	=>	65530,
		16565	=>	65530,
		16566	=>	65530,
		16567	=>	65530,
		16568	=>	65530,
		16569	=>	65530,
		16570	=>	65530,
		16571	=>	65530,
		16572	=>	65530,
		16573	=>	65530,
		16574	=>	65530,
		16575	=>	65530,
		16576	=>	65529,
		16577	=>	65529,
		16578	=>	65529,
		16579	=>	65529,
		16580	=>	65529,
		16581	=>	65529,
		16582	=>	65529,
		16583	=>	65529,
		16584	=>	65529,
		16585	=>	65529,
		16586	=>	65529,
		16587	=>	65529,
		16588	=>	65529,
		16589	=>	65529,
		16590	=>	65529,
		16591	=>	65529,
		16592	=>	65528,
		16593	=>	65528,
		16594	=>	65528,
		16595	=>	65528,
		16596	=>	65528,
		16597	=>	65528,
		16598	=>	65528,
		16599	=>	65528,
		16600	=>	65528,
		16601	=>	65528,
		16602	=>	65528,
		16603	=>	65528,
		16604	=>	65528,
		16605	=>	65528,
		16606	=>	65528,
		16607	=>	65528,
		16608	=>	65527,
		16609	=>	65527,
		16610	=>	65527,
		16611	=>	65527,
		16612	=>	65527,
		16613	=>	65527,
		16614	=>	65527,
		16615	=>	65527,
		16616	=>	65527,
		16617	=>	65527,
		16618	=>	65527,
		16619	=>	65527,
		16620	=>	65527,
		16621	=>	65527,
		16622	=>	65526,
		16623	=>	65526,
		16624	=>	65526,
		16625	=>	65526,
		16626	=>	65526,
		16627	=>	65526,
		16628	=>	65526,
		16629	=>	65526,
		16630	=>	65526,
		16631	=>	65526,
		16632	=>	65526,
		16633	=>	65526,
		16634	=>	65526,
		16635	=>	65526,
		16636	=>	65525,
		16637	=>	65525,
		16638	=>	65525,
		16639	=>	65525,
		16640	=>	65525,
		16641	=>	65525,
		16642	=>	65525,
		16643	=>	65525,
		16644	=>	65525,
		16645	=>	65525,
		16646	=>	65525,
		16647	=>	65525,
		16648	=>	65525,
		16649	=>	65524,
		16650	=>	65524,
		16651	=>	65524,
		16652	=>	65524,
		16653	=>	65524,
		16654	=>	65524,
		16655	=>	65524,
		16656	=>	65524,
		16657	=>	65524,
		16658	=>	65524,
		16659	=>	65524,
		16660	=>	65524,
		16661	=>	65523,
		16662	=>	65523,
		16663	=>	65523,
		16664	=>	65523,
		16665	=>	65523,
		16666	=>	65523,
		16667	=>	65523,
		16668	=>	65523,
		16669	=>	65523,
		16670	=>	65523,
		16671	=>	65523,
		16672	=>	65523,
		16673	=>	65522,
		16674	=>	65522,
		16675	=>	65522,
		16676	=>	65522,
		16677	=>	65522,
		16678	=>	65522,
		16679	=>	65522,
		16680	=>	65522,
		16681	=>	65522,
		16682	=>	65522,
		16683	=>	65522,
		16684	=>	65521,
		16685	=>	65521,
		16686	=>	65521,
		16687	=>	65521,
		16688	=>	65521,
		16689	=>	65521,
		16690	=>	65521,
		16691	=>	65521,
		16692	=>	65521,
		16693	=>	65521,
		16694	=>	65521,
		16695	=>	65520,
		16696	=>	65520,
		16697	=>	65520,
		16698	=>	65520,
		16699	=>	65520,
		16700	=>	65520,
		16701	=>	65520,
		16702	=>	65520,
		16703	=>	65520,
		16704	=>	65520,
		16705	=>	65519,
		16706	=>	65519,
		16707	=>	65519,
		16708	=>	65519,
		16709	=>	65519,
		16710	=>	65519,
		16711	=>	65519,
		16712	=>	65519,
		16713	=>	65519,
		16714	=>	65519,
		16715	=>	65519,
		16716	=>	65518,
		16717	=>	65518,
		16718	=>	65518,
		16719	=>	65518,
		16720	=>	65518,
		16721	=>	65518,
		16722	=>	65518,
		16723	=>	65518,
		16724	=>	65518,
		16725	=>	65517,
		16726	=>	65517,
		16727	=>	65517,
		16728	=>	65517,
		16729	=>	65517,
		16730	=>	65517,
		16731	=>	65517,
		16732	=>	65517,
		16733	=>	65517,
		16734	=>	65517,
		16735	=>	65516,
		16736	=>	65516,
		16737	=>	65516,
		16738	=>	65516,
		16739	=>	65516,
		16740	=>	65516,
		16741	=>	65516,
		16742	=>	65516,
		16743	=>	65516,
		16744	=>	65515,
		16745	=>	65515,
		16746	=>	65515,
		16747	=>	65515,
		16748	=>	65515,
		16749	=>	65515,
		16750	=>	65515,
		16751	=>	65515,
		16752	=>	65515,
		16753	=>	65514,
		16754	=>	65514,
		16755	=>	65514,
		16756	=>	65514,
		16757	=>	65514,
		16758	=>	65514,
		16759	=>	65514,
		16760	=>	65514,
		16761	=>	65514,
		16762	=>	65513,
		16763	=>	65513,
		16764	=>	65513,
		16765	=>	65513,
		16766	=>	65513,
		16767	=>	65513,
		16768	=>	65513,
		16769	=>	65513,
		16770	=>	65513,
		16771	=>	65512,
		16772	=>	65512,
		16773	=>	65512,
		16774	=>	65512,
		16775	=>	65512,
		16776	=>	65512,
		16777	=>	65512,
		16778	=>	65512,
		16779	=>	65512,
		16780	=>	65511,
		16781	=>	65511,
		16782	=>	65511,
		16783	=>	65511,
		16784	=>	65511,
		16785	=>	65511,
		16786	=>	65511,
		16787	=>	65511,
		16788	=>	65510,
		16789	=>	65510,
		16790	=>	65510,
		16791	=>	65510,
		16792	=>	65510,
		16793	=>	65510,
		16794	=>	65510,
		16795	=>	65510,
		16796	=>	65509,
		16797	=>	65509,
		16798	=>	65509,
		16799	=>	65509,
		16800	=>	65509,
		16801	=>	65509,
		16802	=>	65509,
		16803	=>	65509,
		16804	=>	65508,
		16805	=>	65508,
		16806	=>	65508,
		16807	=>	65508,
		16808	=>	65508,
		16809	=>	65508,
		16810	=>	65508,
		16811	=>	65508,
		16812	=>	65507,
		16813	=>	65507,
		16814	=>	65507,
		16815	=>	65507,
		16816	=>	65507,
		16817	=>	65507,
		16818	=>	65507,
		16819	=>	65507,
		16820	=>	65506,
		16821	=>	65506,
		16822	=>	65506,
		16823	=>	65506,
		16824	=>	65506,
		16825	=>	65506,
		16826	=>	65506,
		16827	=>	65505,
		16828	=>	65505,
		16829	=>	65505,
		16830	=>	65505,
		16831	=>	65505,
		16832	=>	65505,
		16833	=>	65505,
		16834	=>	65505,
		16835	=>	65504,
		16836	=>	65504,
		16837	=>	65504,
		16838	=>	65504,
		16839	=>	65504,
		16840	=>	65504,
		16841	=>	65504,
		16842	=>	65503,
		16843	=>	65503,
		16844	=>	65503,
		16845	=>	65503,
		16846	=>	65503,
		16847	=>	65503,
		16848	=>	65503,
		16849	=>	65502,
		16850	=>	65502,
		16851	=>	65502,
		16852	=>	65502,
		16853	=>	65502,
		16854	=>	65502,
		16855	=>	65502,
		16856	=>	65501,
		16857	=>	65501,
		16858	=>	65501,
		16859	=>	65501,
		16860	=>	65501,
		16861	=>	65501,
		16862	=>	65501,
		16863	=>	65500,
		16864	=>	65500,
		16865	=>	65500,
		16866	=>	65500,
		16867	=>	65500,
		16868	=>	65500,
		16869	=>	65500,
		16870	=>	65499,
		16871	=>	65499,
		16872	=>	65499,
		16873	=>	65499,
		16874	=>	65499,
		16875	=>	65499,
		16876	=>	65499,
		16877	=>	65498,
		16878	=>	65498,
		16879	=>	65498,
		16880	=>	65498,
		16881	=>	65498,
		16882	=>	65498,
		16883	=>	65498,
		16884	=>	65497,
		16885	=>	65497,
		16886	=>	65497,
		16887	=>	65497,
		16888	=>	65497,
		16889	=>	65497,
		16890	=>	65496,
		16891	=>	65496,
		16892	=>	65496,
		16893	=>	65496,
		16894	=>	65496,
		16895	=>	65496,
		16896	=>	65496,
		16897	=>	65495,
		16898	=>	65495,
		16899	=>	65495,
		16900	=>	65495,
		16901	=>	65495,
		16902	=>	65495,
		16903	=>	65494,
		16904	=>	65494,
		16905	=>	65494,
		16906	=>	65494,
		16907	=>	65494,
		16908	=>	65494,
		16909	=>	65494,
		16910	=>	65493,
		16911	=>	65493,
		16912	=>	65493,
		16913	=>	65493,
		16914	=>	65493,
		16915	=>	65493,
		16916	=>	65492,
		16917	=>	65492,
		16918	=>	65492,
		16919	=>	65492,
		16920	=>	65492,
		16921	=>	65492,
		16922	=>	65491,
		16923	=>	65491,
		16924	=>	65491,
		16925	=>	65491,
		16926	=>	65491,
		16927	=>	65491,
		16928	=>	65490,
		16929	=>	65490,
		16930	=>	65490,
		16931	=>	65490,
		16932	=>	65490,
		16933	=>	65490,
		16934	=>	65489,
		16935	=>	65489,
		16936	=>	65489,
		16937	=>	65489,
		16938	=>	65489,
		16939	=>	65489,
		16940	=>	65488,
		16941	=>	65488,
		16942	=>	65488,
		16943	=>	65488,
		16944	=>	65488,
		16945	=>	65488,
		16946	=>	65487,
		16947	=>	65487,
		16948	=>	65487,
		16949	=>	65487,
		16950	=>	65487,
		16951	=>	65487,
		16952	=>	65486,
		16953	=>	65486,
		16954	=>	65486,
		16955	=>	65486,
		16956	=>	65486,
		16957	=>	65486,
		16958	=>	65485,
		16959	=>	65485,
		16960	=>	65485,
		16961	=>	65485,
		16962	=>	65485,
		16963	=>	65485,
		16964	=>	65484,
		16965	=>	65484,
		16966	=>	65484,
		16967	=>	65484,
		16968	=>	65484,
		16969	=>	65483,
		16970	=>	65483,
		16971	=>	65483,
		16972	=>	65483,
		16973	=>	65483,
		16974	=>	65483,
		16975	=>	65482,
		16976	=>	65482,
		16977	=>	65482,
		16978	=>	65482,
		16979	=>	65482,
		16980	=>	65482,
		16981	=>	65481,
		16982	=>	65481,
		16983	=>	65481,
		16984	=>	65481,
		16985	=>	65481,
		16986	=>	65480,
		16987	=>	65480,
		16988	=>	65480,
		16989	=>	65480,
		16990	=>	65480,
		16991	=>	65480,
		16992	=>	65479,
		16993	=>	65479,
		16994	=>	65479,
		16995	=>	65479,
		16996	=>	65479,
		16997	=>	65478,
		16998	=>	65478,
		16999	=>	65478,
		17000	=>	65478,
		17001	=>	65478,
		17002	=>	65478,
		17003	=>	65477,
		17004	=>	65477,
		17005	=>	65477,
		17006	=>	65477,
		17007	=>	65477,
		17008	=>	65476,
		17009	=>	65476,
		17010	=>	65476,
		17011	=>	65476,
		17012	=>	65476,
		17013	=>	65475,
		17014	=>	65475,
		17015	=>	65475,
		17016	=>	65475,
		17017	=>	65475,
		17018	=>	65474,
		17019	=>	65474,
		17020	=>	65474,
		17021	=>	65474,
		17022	=>	65474,
		17023	=>	65474,
		17024	=>	65473,
		17025	=>	65473,
		17026	=>	65473,
		17027	=>	65473,
		17028	=>	65473,
		17029	=>	65472,
		17030	=>	65472,
		17031	=>	65472,
		17032	=>	65472,
		17033	=>	65472,
		17034	=>	65471,
		17035	=>	65471,
		17036	=>	65471,
		17037	=>	65471,
		17038	=>	65471,
		17039	=>	65470,
		17040	=>	65470,
		17041	=>	65470,
		17042	=>	65470,
		17043	=>	65470,
		17044	=>	65469,
		17045	=>	65469,
		17046	=>	65469,
		17047	=>	65469,
		17048	=>	65469,
		17049	=>	65468,
		17050	=>	65468,
		17051	=>	65468,
		17052	=>	65468,
		17053	=>	65468,
		17054	=>	65467,
		17055	=>	65467,
		17056	=>	65467,
		17057	=>	65467,
		17058	=>	65467,
		17059	=>	65466,
		17060	=>	65466,
		17061	=>	65466,
		17062	=>	65466,
		17063	=>	65466,
		17064	=>	65465,
		17065	=>	65465,
		17066	=>	65465,
		17067	=>	65465,
		17068	=>	65465,
		17069	=>	65464,
		17070	=>	65464,
		17071	=>	65464,
		17072	=>	65464,
		17073	=>	65464,
		17074	=>	65463,
		17075	=>	65463,
		17076	=>	65463,
		17077	=>	65463,
		17078	=>	65462,
		17079	=>	65462,
		17080	=>	65462,
		17081	=>	65462,
		17082	=>	65462,
		17083	=>	65461,
		17084	=>	65461,
		17085	=>	65461,
		17086	=>	65461,
		17087	=>	65461,
		17088	=>	65460,
		17089	=>	65460,
		17090	=>	65460,
		17091	=>	65460,
		17092	=>	65460,
		17093	=>	65459,
		17094	=>	65459,
		17095	=>	65459,
		17096	=>	65459,
		17097	=>	65458,
		17098	=>	65458,
		17099	=>	65458,
		17100	=>	65458,
		17101	=>	65458,
		17102	=>	65457,
		17103	=>	65457,
		17104	=>	65457,
		17105	=>	65457,
		17106	=>	65457,
		17107	=>	65456,
		17108	=>	65456,
		17109	=>	65456,
		17110	=>	65456,
		17111	=>	65455,
		17112	=>	65455,
		17113	=>	65455,
		17114	=>	65455,
		17115	=>	65455,
		17116	=>	65454,
		17117	=>	65454,
		17118	=>	65454,
		17119	=>	65454,
		17120	=>	65453,
		17121	=>	65453,
		17122	=>	65453,
		17123	=>	65453,
		17124	=>	65453,
		17125	=>	65452,
		17126	=>	65452,
		17127	=>	65452,
		17128	=>	65452,
		17129	=>	65451,
		17130	=>	65451,
		17131	=>	65451,
		17132	=>	65451,
		17133	=>	65451,
		17134	=>	65450,
		17135	=>	65450,
		17136	=>	65450,
		17137	=>	65450,
		17138	=>	65449,
		17139	=>	65449,
		17140	=>	65449,
		17141	=>	65449,
		17142	=>	65449,
		17143	=>	65448,
		17144	=>	65448,
		17145	=>	65448,
		17146	=>	65448,
		17147	=>	65447,
		17148	=>	65447,
		17149	=>	65447,
		17150	=>	65447,
		17151	=>	65446,
		17152	=>	65446,
		17153	=>	65446,
		17154	=>	65446,
		17155	=>	65446,
		17156	=>	65445,
		17157	=>	65445,
		17158	=>	65445,
		17159	=>	65445,
		17160	=>	65444,
		17161	=>	65444,
		17162	=>	65444,
		17163	=>	65444,
		17164	=>	65443,
		17165	=>	65443,
		17166	=>	65443,
		17167	=>	65443,
		17168	=>	65442,
		17169	=>	65442,
		17170	=>	65442,
		17171	=>	65442,
		17172	=>	65442,
		17173	=>	65441,
		17174	=>	65441,
		17175	=>	65441,
		17176	=>	65441,
		17177	=>	65440,
		17178	=>	65440,
		17179	=>	65440,
		17180	=>	65440,
		17181	=>	65439,
		17182	=>	65439,
		17183	=>	65439,
		17184	=>	65439,
		17185	=>	65438,
		17186	=>	65438,
		17187	=>	65438,
		17188	=>	65438,
		17189	=>	65437,
		17190	=>	65437,
		17191	=>	65437,
		17192	=>	65437,
		17193	=>	65436,
		17194	=>	65436,
		17195	=>	65436,
		17196	=>	65436,
		17197	=>	65436,
		17198	=>	65435,
		17199	=>	65435,
		17200	=>	65435,
		17201	=>	65435,
		17202	=>	65434,
		17203	=>	65434,
		17204	=>	65434,
		17205	=>	65434,
		17206	=>	65433,
		17207	=>	65433,
		17208	=>	65433,
		17209	=>	65433,
		17210	=>	65432,
		17211	=>	65432,
		17212	=>	65432,
		17213	=>	65432,
		17214	=>	65431,
		17215	=>	65431,
		17216	=>	65431,
		17217	=>	65431,
		17218	=>	65430,
		17219	=>	65430,
		17220	=>	65430,
		17221	=>	65430,
		17222	=>	65429,
		17223	=>	65429,
		17224	=>	65429,
		17225	=>	65429,
		17226	=>	65428,
		17227	=>	65428,
		17228	=>	65428,
		17229	=>	65428,
		17230	=>	65427,
		17231	=>	65427,
		17232	=>	65427,
		17233	=>	65427,
		17234	=>	65426,
		17235	=>	65426,
		17236	=>	65426,
		17237	=>	65425,
		17238	=>	65425,
		17239	=>	65425,
		17240	=>	65425,
		17241	=>	65424,
		17242	=>	65424,
		17243	=>	65424,
		17244	=>	65424,
		17245	=>	65423,
		17246	=>	65423,
		17247	=>	65423,
		17248	=>	65423,
		17249	=>	65422,
		17250	=>	65422,
		17251	=>	65422,
		17252	=>	65422,
		17253	=>	65421,
		17254	=>	65421,
		17255	=>	65421,
		17256	=>	65421,
		17257	=>	65420,
		17258	=>	65420,
		17259	=>	65420,
		17260	=>	65420,
		17261	=>	65419,
		17262	=>	65419,
		17263	=>	65419,
		17264	=>	65418,
		17265	=>	65418,
		17266	=>	65418,
		17267	=>	65418,
		17268	=>	65417,
		17269	=>	65417,
		17270	=>	65417,
		17271	=>	65417,
		17272	=>	65416,
		17273	=>	65416,
		17274	=>	65416,
		17275	=>	65416,
		17276	=>	65415,
		17277	=>	65415,
		17278	=>	65415,
		17279	=>	65414,
		17280	=>	65414,
		17281	=>	65414,
		17282	=>	65414,
		17283	=>	65413,
		17284	=>	65413,
		17285	=>	65413,
		17286	=>	65413,
		17287	=>	65412,
		17288	=>	65412,
		17289	=>	65412,
		17290	=>	65411,
		17291	=>	65411,
		17292	=>	65411,
		17293	=>	65411,
		17294	=>	65410,
		17295	=>	65410,
		17296	=>	65410,
		17297	=>	65410,
		17298	=>	65409,
		17299	=>	65409,
		17300	=>	65409,
		17301	=>	65408,
		17302	=>	65408,
		17303	=>	65408,
		17304	=>	65408,
		17305	=>	65407,
		17306	=>	65407,
		17307	=>	65407,
		17308	=>	65407,
		17309	=>	65406,
		17310	=>	65406,
		17311	=>	65406,
		17312	=>	65405,
		17313	=>	65405,
		17314	=>	65405,
		17315	=>	65405,
		17316	=>	65404,
		17317	=>	65404,
		17318	=>	65404,
		17319	=>	65403,
		17320	=>	65403,
		17321	=>	65403,
		17322	=>	65403,
		17323	=>	65402,
		17324	=>	65402,
		17325	=>	65402,
		17326	=>	65401,
		17327	=>	65401,
		17328	=>	65401,
		17329	=>	65401,
		17330	=>	65400,
		17331	=>	65400,
		17332	=>	65400,
		17333	=>	65399,
		17334	=>	65399,
		17335	=>	65399,
		17336	=>	65399,
		17337	=>	65398,
		17338	=>	65398,
		17339	=>	65398,
		17340	=>	65397,
		17341	=>	65397,
		17342	=>	65397,
		17343	=>	65397,
		17344	=>	65396,
		17345	=>	65396,
		17346	=>	65396,
		17347	=>	65395,
		17348	=>	65395,
		17349	=>	65395,
		17350	=>	65395,
		17351	=>	65394,
		17352	=>	65394,
		17353	=>	65394,
		17354	=>	65393,
		17355	=>	65393,
		17356	=>	65393,
		17357	=>	65393,
		17358	=>	65392,
		17359	=>	65392,
		17360	=>	65392,
		17361	=>	65391,
		17362	=>	65391,
		17363	=>	65391,
		17364	=>	65390,
		17365	=>	65390,
		17366	=>	65390,
		17367	=>	65390,
		17368	=>	65389,
		17369	=>	65389,
		17370	=>	65389,
		17371	=>	65388,
		17372	=>	65388,
		17373	=>	65388,
		17374	=>	65388,
		17375	=>	65387,
		17376	=>	65387,
		17377	=>	65387,
		17378	=>	65386,
		17379	=>	65386,
		17380	=>	65386,
		17381	=>	65385,
		17382	=>	65385,
		17383	=>	65385,
		17384	=>	65385,
		17385	=>	65384,
		17386	=>	65384,
		17387	=>	65384,
		17388	=>	65383,
		17389	=>	65383,
		17390	=>	65383,
		17391	=>	65382,
		17392	=>	65382,
		17393	=>	65382,
		17394	=>	65381,
		17395	=>	65381,
		17396	=>	65381,
		17397	=>	65381,
		17398	=>	65380,
		17399	=>	65380,
		17400	=>	65380,
		17401	=>	65379,
		17402	=>	65379,
		17403	=>	65379,
		17404	=>	65378,
		17405	=>	65378,
		17406	=>	65378,
		17407	=>	65378,
		17408	=>	65377,
		17409	=>	65377,
		17410	=>	65377,
		17411	=>	65376,
		17412	=>	65376,
		17413	=>	65376,
		17414	=>	65375,
		17415	=>	65375,
		17416	=>	65375,
		17417	=>	65374,
		17418	=>	65374,
		17419	=>	65374,
		17420	=>	65373,
		17421	=>	65373,
		17422	=>	65373,
		17423	=>	65373,
		17424	=>	65372,
		17425	=>	65372,
		17426	=>	65372,
		17427	=>	65371,
		17428	=>	65371,
		17429	=>	65371,
		17430	=>	65370,
		17431	=>	65370,
		17432	=>	65370,
		17433	=>	65369,
		17434	=>	65369,
		17435	=>	65369,
		17436	=>	65368,
		17437	=>	65368,
		17438	=>	65368,
		17439	=>	65368,
		17440	=>	65367,
		17441	=>	65367,
		17442	=>	65367,
		17443	=>	65366,
		17444	=>	65366,
		17445	=>	65366,
		17446	=>	65365,
		17447	=>	65365,
		17448	=>	65365,
		17449	=>	65364,
		17450	=>	65364,
		17451	=>	65364,
		17452	=>	65363,
		17453	=>	65363,
		17454	=>	65363,
		17455	=>	65362,
		17456	=>	65362,
		17457	=>	65362,
		17458	=>	65361,
		17459	=>	65361,
		17460	=>	65361,
		17461	=>	65360,
		17462	=>	65360,
		17463	=>	65360,
		17464	=>	65360,
		17465	=>	65359,
		17466	=>	65359,
		17467	=>	65359,
		17468	=>	65358,
		17469	=>	65358,
		17470	=>	65358,
		17471	=>	65357,
		17472	=>	65357,
		17473	=>	65357,
		17474	=>	65356,
		17475	=>	65356,
		17476	=>	65356,
		17477	=>	65355,
		17478	=>	65355,
		17479	=>	65355,
		17480	=>	65354,
		17481	=>	65354,
		17482	=>	65354,
		17483	=>	65353,
		17484	=>	65353,
		17485	=>	65353,
		17486	=>	65352,
		17487	=>	65352,
		17488	=>	65352,
		17489	=>	65351,
		17490	=>	65351,
		17491	=>	65351,
		17492	=>	65350,
		17493	=>	65350,
		17494	=>	65350,
		17495	=>	65349,
		17496	=>	65349,
		17497	=>	65349,
		17498	=>	65348,
		17499	=>	65348,
		17500	=>	65348,
		17501	=>	65347,
		17502	=>	65347,
		17503	=>	65347,
		17504	=>	65346,
		17505	=>	65346,
		17506	=>	65346,
		17507	=>	65345,
		17508	=>	65345,
		17509	=>	65345,
		17510	=>	65344,
		17511	=>	65344,
		17512	=>	65344,
		17513	=>	65343,
		17514	=>	65343,
		17515	=>	65343,
		17516	=>	65342,
		17517	=>	65342,
		17518	=>	65342,
		17519	=>	65341,
		17520	=>	65341,
		17521	=>	65341,
		17522	=>	65340,
		17523	=>	65340,
		17524	=>	65339,
		17525	=>	65339,
		17526	=>	65339,
		17527	=>	65338,
		17528	=>	65338,
		17529	=>	65338,
		17530	=>	65337,
		17531	=>	65337,
		17532	=>	65337,
		17533	=>	65336,
		17534	=>	65336,
		17535	=>	65336,
		17536	=>	65335,
		17537	=>	65335,
		17538	=>	65335,
		17539	=>	65334,
		17540	=>	65334,
		17541	=>	65334,
		17542	=>	65333,
		17543	=>	65333,
		17544	=>	65333,
		17545	=>	65332,
		17546	=>	65332,
		17547	=>	65332,
		17548	=>	65331,
		17549	=>	65331,
		17550	=>	65330,
		17551	=>	65330,
		17552	=>	65330,
		17553	=>	65329,
		17554	=>	65329,
		17555	=>	65329,
		17556	=>	65328,
		17557	=>	65328,
		17558	=>	65328,
		17559	=>	65327,
		17560	=>	65327,
		17561	=>	65327,
		17562	=>	65326,
		17563	=>	65326,
		17564	=>	65326,
		17565	=>	65325,
		17566	=>	65325,
		17567	=>	65324,
		17568	=>	65324,
		17569	=>	65324,
		17570	=>	65323,
		17571	=>	65323,
		17572	=>	65323,
		17573	=>	65322,
		17574	=>	65322,
		17575	=>	65322,
		17576	=>	65321,
		17577	=>	65321,
		17578	=>	65321,
		17579	=>	65320,
		17580	=>	65320,
		17581	=>	65319,
		17582	=>	65319,
		17583	=>	65319,
		17584	=>	65318,
		17585	=>	65318,
		17586	=>	65318,
		17587	=>	65317,
		17588	=>	65317,
		17589	=>	65317,
		17590	=>	65316,
		17591	=>	65316,
		17592	=>	65315,
		17593	=>	65315,
		17594	=>	65315,
		17595	=>	65314,
		17596	=>	65314,
		17597	=>	65314,
		17598	=>	65313,
		17599	=>	65313,
		17600	=>	65313,
		17601	=>	65312,
		17602	=>	65312,
		17603	=>	65311,
		17604	=>	65311,
		17605	=>	65311,
		17606	=>	65310,
		17607	=>	65310,
		17608	=>	65310,
		17609	=>	65309,
		17610	=>	65309,
		17611	=>	65309,
		17612	=>	65308,
		17613	=>	65308,
		17614	=>	65307,
		17615	=>	65307,
		17616	=>	65307,
		17617	=>	65306,
		17618	=>	65306,
		17619	=>	65306,
		17620	=>	65305,
		17621	=>	65305,
		17622	=>	65304,
		17623	=>	65304,
		17624	=>	65304,
		17625	=>	65303,
		17626	=>	65303,
		17627	=>	65303,
		17628	=>	65302,
		17629	=>	65302,
		17630	=>	65301,
		17631	=>	65301,
		17632	=>	65301,
		17633	=>	65300,
		17634	=>	65300,
		17635	=>	65300,
		17636	=>	65299,
		17637	=>	65299,
		17638	=>	65298,
		17639	=>	65298,
		17640	=>	65298,
		17641	=>	65297,
		17642	=>	65297,
		17643	=>	65297,
		17644	=>	65296,
		17645	=>	65296,
		17646	=>	65295,
		17647	=>	65295,
		17648	=>	65295,
		17649	=>	65294,
		17650	=>	65294,
		17651	=>	65294,
		17652	=>	65293,
		17653	=>	65293,
		17654	=>	65292,
		17655	=>	65292,
		17656	=>	65292,
		17657	=>	65291,
		17658	=>	65291,
		17659	=>	65290,
		17660	=>	65290,
		17661	=>	65290,
		17662	=>	65289,
		17663	=>	65289,
		17664	=>	65289,
		17665	=>	65288,
		17666	=>	65288,
		17667	=>	65287,
		17668	=>	65287,
		17669	=>	65287,
		17670	=>	65286,
		17671	=>	65286,
		17672	=>	65285,
		17673	=>	65285,
		17674	=>	65285,
		17675	=>	65284,
		17676	=>	65284,
		17677	=>	65284,
		17678	=>	65283,
		17679	=>	65283,
		17680	=>	65282,
		17681	=>	65282,
		17682	=>	65282,
		17683	=>	65281,
		17684	=>	65281,
		17685	=>	65280,
		17686	=>	65280,
		17687	=>	65280,
		17688	=>	65279,
		17689	=>	65279,
		17690	=>	65278,
		17691	=>	65278,
		17692	=>	65278,
		17693	=>	65277,
		17694	=>	65277,
		17695	=>	65277,
		17696	=>	65276,
		17697	=>	65276,
		17698	=>	65275,
		17699	=>	65275,
		17700	=>	65275,
		17701	=>	65274,
		17702	=>	65274,
		17703	=>	65273,
		17704	=>	65273,
		17705	=>	65273,
		17706	=>	65272,
		17707	=>	65272,
		17708	=>	65271,
		17709	=>	65271,
		17710	=>	65271,
		17711	=>	65270,
		17712	=>	65270,
		17713	=>	65269,
		17714	=>	65269,
		17715	=>	65269,
		17716	=>	65268,
		17717	=>	65268,
		17718	=>	65267,
		17719	=>	65267,
		17720	=>	65267,
		17721	=>	65266,
		17722	=>	65266,
		17723	=>	65265,
		17724	=>	65265,
		17725	=>	65265,
		17726	=>	65264,
		17727	=>	65264,
		17728	=>	65263,
		17729	=>	65263,
		17730	=>	65263,
		17731	=>	65262,
		17732	=>	65262,
		17733	=>	65261,
		17734	=>	65261,
		17735	=>	65261,
		17736	=>	65260,
		17737	=>	65260,
		17738	=>	65259,
		17739	=>	65259,
		17740	=>	65258,
		17741	=>	65258,
		17742	=>	65258,
		17743	=>	65257,
		17744	=>	65257,
		17745	=>	65256,
		17746	=>	65256,
		17747	=>	65256,
		17748	=>	65255,
		17749	=>	65255,
		17750	=>	65254,
		17751	=>	65254,
		17752	=>	65254,
		17753	=>	65253,
		17754	=>	65253,
		17755	=>	65252,
		17756	=>	65252,
		17757	=>	65252,
		17758	=>	65251,
		17759	=>	65251,
		17760	=>	65250,
		17761	=>	65250,
		17762	=>	65249,
		17763	=>	65249,
		17764	=>	65249,
		17765	=>	65248,
		17766	=>	65248,
		17767	=>	65247,
		17768	=>	65247,
		17769	=>	65247,
		17770	=>	65246,
		17771	=>	65246,
		17772	=>	65245,
		17773	=>	65245,
		17774	=>	65244,
		17775	=>	65244,
		17776	=>	65244,
		17777	=>	65243,
		17778	=>	65243,
		17779	=>	65242,
		17780	=>	65242,
		17781	=>	65242,
		17782	=>	65241,
		17783	=>	65241,
		17784	=>	65240,
		17785	=>	65240,
		17786	=>	65239,
		17787	=>	65239,
		17788	=>	65239,
		17789	=>	65238,
		17790	=>	65238,
		17791	=>	65237,
		17792	=>	65237,
		17793	=>	65236,
		17794	=>	65236,
		17795	=>	65236,
		17796	=>	65235,
		17797	=>	65235,
		17798	=>	65234,
		17799	=>	65234,
		17800	=>	65234,
		17801	=>	65233,
		17802	=>	65233,
		17803	=>	65232,
		17804	=>	65232,
		17805	=>	65231,
		17806	=>	65231,
		17807	=>	65231,
		17808	=>	65230,
		17809	=>	65230,
		17810	=>	65229,
		17811	=>	65229,
		17812	=>	65228,
		17813	=>	65228,
		17814	=>	65228,
		17815	=>	65227,
		17816	=>	65227,
		17817	=>	65226,
		17818	=>	65226,
		17819	=>	65225,
		17820	=>	65225,
		17821	=>	65225,
		17822	=>	65224,
		17823	=>	65224,
		17824	=>	65223,
		17825	=>	65223,
		17826	=>	65222,
		17827	=>	65222,
		17828	=>	65221,
		17829	=>	65221,
		17830	=>	65221,
		17831	=>	65220,
		17832	=>	65220,
		17833	=>	65219,
		17834	=>	65219,
		17835	=>	65218,
		17836	=>	65218,
		17837	=>	65218,
		17838	=>	65217,
		17839	=>	65217,
		17840	=>	65216,
		17841	=>	65216,
		17842	=>	65215,
		17843	=>	65215,
		17844	=>	65215,
		17845	=>	65214,
		17846	=>	65214,
		17847	=>	65213,
		17848	=>	65213,
		17849	=>	65212,
		17850	=>	65212,
		17851	=>	65211,
		17852	=>	65211,
		17853	=>	65211,
		17854	=>	65210,
		17855	=>	65210,
		17856	=>	65209,
		17857	=>	65209,
		17858	=>	65208,
		17859	=>	65208,
		17860	=>	65207,
		17861	=>	65207,
		17862	=>	65207,
		17863	=>	65206,
		17864	=>	65206,
		17865	=>	65205,
		17866	=>	65205,
		17867	=>	65204,
		17868	=>	65204,
		17869	=>	65203,
		17870	=>	65203,
		17871	=>	65203,
		17872	=>	65202,
		17873	=>	65202,
		17874	=>	65201,
		17875	=>	65201,
		17876	=>	65200,
		17877	=>	65200,
		17878	=>	65199,
		17879	=>	65199,
		17880	=>	65199,
		17881	=>	65198,
		17882	=>	65198,
		17883	=>	65197,
		17884	=>	65197,
		17885	=>	65196,
		17886	=>	65196,
		17887	=>	65195,
		17888	=>	65195,
		17889	=>	65194,
		17890	=>	65194,
		17891	=>	65194,
		17892	=>	65193,
		17893	=>	65193,
		17894	=>	65192,
		17895	=>	65192,
		17896	=>	65191,
		17897	=>	65191,
		17898	=>	65190,
		17899	=>	65190,
		17900	=>	65190,
		17901	=>	65189,
		17902	=>	65189,
		17903	=>	65188,
		17904	=>	65188,
		17905	=>	65187,
		17906	=>	65187,
		17907	=>	65186,
		17908	=>	65186,
		17909	=>	65185,
		17910	=>	65185,
		17911	=>	65184,
		17912	=>	65184,
		17913	=>	65184,
		17914	=>	65183,
		17915	=>	65183,
		17916	=>	65182,
		17917	=>	65182,
		17918	=>	65181,
		17919	=>	65181,
		17920	=>	65180,
		17921	=>	65180,
		17922	=>	65179,
		17923	=>	65179,
		17924	=>	65178,
		17925	=>	65178,
		17926	=>	65178,
		17927	=>	65177,
		17928	=>	65177,
		17929	=>	65176,
		17930	=>	65176,
		17931	=>	65175,
		17932	=>	65175,
		17933	=>	65174,
		17934	=>	65174,
		17935	=>	65173,
		17936	=>	65173,
		17937	=>	65172,
		17938	=>	65172,
		17939	=>	65172,
		17940	=>	65171,
		17941	=>	65171,
		17942	=>	65170,
		17943	=>	65170,
		17944	=>	65169,
		17945	=>	65169,
		17946	=>	65168,
		17947	=>	65168,
		17948	=>	65167,
		17949	=>	65167,
		17950	=>	65166,
		17951	=>	65166,
		17952	=>	65165,
		17953	=>	65165,
		17954	=>	65164,
		17955	=>	65164,
		17956	=>	65164,
		17957	=>	65163,
		17958	=>	65163,
		17959	=>	65162,
		17960	=>	65162,
		17961	=>	65161,
		17962	=>	65161,
		17963	=>	65160,
		17964	=>	65160,
		17965	=>	65159,
		17966	=>	65159,
		17967	=>	65158,
		17968	=>	65158,
		17969	=>	65157,
		17970	=>	65157,
		17971	=>	65156,
		17972	=>	65156,
		17973	=>	65155,
		17974	=>	65155,
		17975	=>	65155,
		17976	=>	65154,
		17977	=>	65154,
		17978	=>	65153,
		17979	=>	65153,
		17980	=>	65152,
		17981	=>	65152,
		17982	=>	65151,
		17983	=>	65151,
		17984	=>	65150,
		17985	=>	65150,
		17986	=>	65149,
		17987	=>	65149,
		17988	=>	65148,
		17989	=>	65148,
		17990	=>	65147,
		17991	=>	65147,
		17992	=>	65146,
		17993	=>	65146,
		17994	=>	65145,
		17995	=>	65145,
		17996	=>	65144,
		17997	=>	65144,
		17998	=>	65143,
		17999	=>	65143,
		18000	=>	65143,
		18001	=>	65142,
		18002	=>	65142,
		18003	=>	65141,
		18004	=>	65141,
		18005	=>	65140,
		18006	=>	65140,
		18007	=>	65139,
		18008	=>	65139,
		18009	=>	65138,
		18010	=>	65138,
		18011	=>	65137,
		18012	=>	65137,
		18013	=>	65136,
		18014	=>	65136,
		18015	=>	65135,
		18016	=>	65135,
		18017	=>	65134,
		18018	=>	65134,
		18019	=>	65133,
		18020	=>	65133,
		18021	=>	65132,
		18022	=>	65132,
		18023	=>	65131,
		18024	=>	65131,
		18025	=>	65130,
		18026	=>	65130,
		18027	=>	65129,
		18028	=>	65129,
		18029	=>	65128,
		18030	=>	65128,
		18031	=>	65127,
		18032	=>	65127,
		18033	=>	65126,
		18034	=>	65126,
		18035	=>	65125,
		18036	=>	65125,
		18037	=>	65124,
		18038	=>	65124,
		18039	=>	65123,
		18040	=>	65123,
		18041	=>	65122,
		18042	=>	65122,
		18043	=>	65121,
		18044	=>	65121,
		18045	=>	65120,
		18046	=>	65120,
		18047	=>	65119,
		18048	=>	65119,
		18049	=>	65118,
		18050	=>	65118,
		18051	=>	65117,
		18052	=>	65117,
		18053	=>	65116,
		18054	=>	65116,
		18055	=>	65115,
		18056	=>	65115,
		18057	=>	65114,
		18058	=>	65114,
		18059	=>	65113,
		18060	=>	65113,
		18061	=>	65112,
		18062	=>	65112,
		18063	=>	65111,
		18064	=>	65111,
		18065	=>	65110,
		18066	=>	65110,
		18067	=>	65109,
		18068	=>	65109,
		18069	=>	65108,
		18070	=>	65108,
		18071	=>	65107,
		18072	=>	65107,
		18073	=>	65106,
		18074	=>	65106,
		18075	=>	65105,
		18076	=>	65105,
		18077	=>	65104,
		18078	=>	65104,
		18079	=>	65103,
		18080	=>	65103,
		18081	=>	65102,
		18082	=>	65102,
		18083	=>	65101,
		18084	=>	65101,
		18085	=>	65100,
		18086	=>	65100,
		18087	=>	65099,
		18088	=>	65099,
		18089	=>	65098,
		18090	=>	65098,
		18091	=>	65097,
		18092	=>	65097,
		18093	=>	65096,
		18094	=>	65096,
		18095	=>	65095,
		18096	=>	65095,
		18097	=>	65094,
		18098	=>	65094,
		18099	=>	65093,
		18100	=>	65093,
		18101	=>	65092,
		18102	=>	65092,
		18103	=>	65091,
		18104	=>	65090,
		18105	=>	65090,
		18106	=>	65089,
		18107	=>	65089,
		18108	=>	65088,
		18109	=>	65088,
		18110	=>	65087,
		18111	=>	65087,
		18112	=>	65086,
		18113	=>	65086,
		18114	=>	65085,
		18115	=>	65085,
		18116	=>	65084,
		18117	=>	65084,
		18118	=>	65083,
		18119	=>	65083,
		18120	=>	65082,
		18121	=>	65082,
		18122	=>	65081,
		18123	=>	65081,
		18124	=>	65080,
		18125	=>	65080,
		18126	=>	65079,
		18127	=>	65079,
		18128	=>	65078,
		18129	=>	65078,
		18130	=>	65077,
		18131	=>	65076,
		18132	=>	65076,
		18133	=>	65075,
		18134	=>	65075,
		18135	=>	65074,
		18136	=>	65074,
		18137	=>	65073,
		18138	=>	65073,
		18139	=>	65072,
		18140	=>	65072,
		18141	=>	65071,
		18142	=>	65071,
		18143	=>	65070,
		18144	=>	65070,
		18145	=>	65069,
		18146	=>	65069,
		18147	=>	65068,
		18148	=>	65068,
		18149	=>	65067,
		18150	=>	65066,
		18151	=>	65066,
		18152	=>	65065,
		18153	=>	65065,
		18154	=>	65064,
		18155	=>	65064,
		18156	=>	65063,
		18157	=>	65063,
		18158	=>	65062,
		18159	=>	65062,
		18160	=>	65061,
		18161	=>	65061,
		18162	=>	65060,
		18163	=>	65060,
		18164	=>	65059,
		18165	=>	65058,
		18166	=>	65058,
		18167	=>	65057,
		18168	=>	65057,
		18169	=>	65056,
		18170	=>	65056,
		18171	=>	65055,
		18172	=>	65055,
		18173	=>	65054,
		18174	=>	65054,
		18175	=>	65053,
		18176	=>	65053,
		18177	=>	65052,
		18178	=>	65052,
		18179	=>	65051,
		18180	=>	65050,
		18181	=>	65050,
		18182	=>	65049,
		18183	=>	65049,
		18184	=>	65048,
		18185	=>	65048,
		18186	=>	65047,
		18187	=>	65047,
		18188	=>	65046,
		18189	=>	65046,
		18190	=>	65045,
		18191	=>	65044,
		18192	=>	65044,
		18193	=>	65043,
		18194	=>	65043,
		18195	=>	65042,
		18196	=>	65042,
		18197	=>	65041,
		18198	=>	65041,
		18199	=>	65040,
		18200	=>	65040,
		18201	=>	65039,
		18202	=>	65039,
		18203	=>	65038,
		18204	=>	65037,
		18205	=>	65037,
		18206	=>	65036,
		18207	=>	65036,
		18208	=>	65035,
		18209	=>	65035,
		18210	=>	65034,
		18211	=>	65034,
		18212	=>	65033,
		18213	=>	65033,
		18214	=>	65032,
		18215	=>	65031,
		18216	=>	65031,
		18217	=>	65030,
		18218	=>	65030,
		18219	=>	65029,
		18220	=>	65029,
		18221	=>	65028,
		18222	=>	65028,
		18223	=>	65027,
		18224	=>	65026,
		18225	=>	65026,
		18226	=>	65025,
		18227	=>	65025,
		18228	=>	65024,
		18229	=>	65024,
		18230	=>	65023,
		18231	=>	65023,
		18232	=>	65022,
		18233	=>	65021,
		18234	=>	65021,
		18235	=>	65020,
		18236	=>	65020,
		18237	=>	65019,
		18238	=>	65019,
		18239	=>	65018,
		18240	=>	65018,
		18241	=>	65017,
		18242	=>	65016,
		18243	=>	65016,
		18244	=>	65015,
		18245	=>	65015,
		18246	=>	65014,
		18247	=>	65014,
		18248	=>	65013,
		18249	=>	65013,
		18250	=>	65012,
		18251	=>	65011,
		18252	=>	65011,
		18253	=>	65010,
		18254	=>	65010,
		18255	=>	65009,
		18256	=>	65009,
		18257	=>	65008,
		18258	=>	65008,
		18259	=>	65007,
		18260	=>	65006,
		18261	=>	65006,
		18262	=>	65005,
		18263	=>	65005,
		18264	=>	65004,
		18265	=>	65004,
		18266	=>	65003,
		18267	=>	65002,
		18268	=>	65002,
		18269	=>	65001,
		18270	=>	65001,
		18271	=>	65000,
		18272	=>	65000,
		18273	=>	64999,
		18274	=>	64999,
		18275	=>	64998,
		18276	=>	64997,
		18277	=>	64997,
		18278	=>	64996,
		18279	=>	64996,
		18280	=>	64995,
		18281	=>	64995,
		18282	=>	64994,
		18283	=>	64993,
		18284	=>	64993,
		18285	=>	64992,
		18286	=>	64992,
		18287	=>	64991,
		18288	=>	64991,
		18289	=>	64990,
		18290	=>	64989,
		18291	=>	64989,
		18292	=>	64988,
		18293	=>	64988,
		18294	=>	64987,
		18295	=>	64987,
		18296	=>	64986,
		18297	=>	64985,
		18298	=>	64985,
		18299	=>	64984,
		18300	=>	64984,
		18301	=>	64983,
		18302	=>	64983,
		18303	=>	64982,
		18304	=>	64981,
		18305	=>	64981,
		18306	=>	64980,
		18307	=>	64980,
		18308	=>	64979,
		18309	=>	64979,
		18310	=>	64978,
		18311	=>	64977,
		18312	=>	64977,
		18313	=>	64976,
		18314	=>	64976,
		18315	=>	64975,
		18316	=>	64974,
		18317	=>	64974,
		18318	=>	64973,
		18319	=>	64973,
		18320	=>	64972,
		18321	=>	64972,
		18322	=>	64971,
		18323	=>	64970,
		18324	=>	64970,
		18325	=>	64969,
		18326	=>	64969,
		18327	=>	64968,
		18328	=>	64968,
		18329	=>	64967,
		18330	=>	64966,
		18331	=>	64966,
		18332	=>	64965,
		18333	=>	64965,
		18334	=>	64964,
		18335	=>	64963,
		18336	=>	64963,
		18337	=>	64962,
		18338	=>	64962,
		18339	=>	64961,
		18340	=>	64961,
		18341	=>	64960,
		18342	=>	64959,
		18343	=>	64959,
		18344	=>	64958,
		18345	=>	64958,
		18346	=>	64957,
		18347	=>	64956,
		18348	=>	64956,
		18349	=>	64955,
		18350	=>	64955,
		18351	=>	64954,
		18352	=>	64953,
		18353	=>	64953,
		18354	=>	64952,
		18355	=>	64952,
		18356	=>	64951,
		18357	=>	64951,
		18358	=>	64950,
		18359	=>	64949,
		18360	=>	64949,
		18361	=>	64948,
		18362	=>	64948,
		18363	=>	64947,
		18364	=>	64946,
		18365	=>	64946,
		18366	=>	64945,
		18367	=>	64945,
		18368	=>	64944,
		18369	=>	64943,
		18370	=>	64943,
		18371	=>	64942,
		18372	=>	64942,
		18373	=>	64941,
		18374	=>	64940,
		18375	=>	64940,
		18376	=>	64939,
		18377	=>	64939,
		18378	=>	64938,
		18379	=>	64937,
		18380	=>	64937,
		18381	=>	64936,
		18382	=>	64936,
		18383	=>	64935,
		18384	=>	64934,
		18385	=>	64934,
		18386	=>	64933,
		18387	=>	64933,
		18388	=>	64932,
		18389	=>	64931,
		18390	=>	64931,
		18391	=>	64930,
		18392	=>	64930,
		18393	=>	64929,
		18394	=>	64928,
		18395	=>	64928,
		18396	=>	64927,
		18397	=>	64927,
		18398	=>	64926,
		18399	=>	64925,
		18400	=>	64925,
		18401	=>	64924,
		18402	=>	64924,
		18403	=>	64923,
		18404	=>	64922,
		18405	=>	64922,
		18406	=>	64921,
		18407	=>	64921,
		18408	=>	64920,
		18409	=>	64919,
		18410	=>	64919,
		18411	=>	64918,
		18412	=>	64918,
		18413	=>	64917,
		18414	=>	64916,
		18415	=>	64916,
		18416	=>	64915,
		18417	=>	64915,
		18418	=>	64914,
		18419	=>	64913,
		18420	=>	64913,
		18421	=>	64912,
		18422	=>	64911,
		18423	=>	64911,
		18424	=>	64910,
		18425	=>	64910,
		18426	=>	64909,
		18427	=>	64908,
		18428	=>	64908,
		18429	=>	64907,
		18430	=>	64907,
		18431	=>	64906,
		18432	=>	64905,
		18433	=>	64905,
		18434	=>	64904,
		18435	=>	64904,
		18436	=>	64903,
		18437	=>	64902,
		18438	=>	64902,
		18439	=>	64901,
		18440	=>	64900,
		18441	=>	64900,
		18442	=>	64899,
		18443	=>	64899,
		18444	=>	64898,
		18445	=>	64897,
		18446	=>	64897,
		18447	=>	64896,
		18448	=>	64896,
		18449	=>	64895,
		18450	=>	64894,
		18451	=>	64894,
		18452	=>	64893,
		18453	=>	64892,
		18454	=>	64892,
		18455	=>	64891,
		18456	=>	64891,
		18457	=>	64890,
		18458	=>	64889,
		18459	=>	64889,
		18460	=>	64888,
		18461	=>	64887,
		18462	=>	64887,
		18463	=>	64886,
		18464	=>	64886,
		18465	=>	64885,
		18466	=>	64884,
		18467	=>	64884,
		18468	=>	64883,
		18469	=>	64883,
		18470	=>	64882,
		18471	=>	64881,
		18472	=>	64881,
		18473	=>	64880,
		18474	=>	64879,
		18475	=>	64879,
		18476	=>	64878,
		18477	=>	64878,
		18478	=>	64877,
		18479	=>	64876,
		18480	=>	64876,
		18481	=>	64875,
		18482	=>	64874,
		18483	=>	64874,
		18484	=>	64873,
		18485	=>	64872,
		18486	=>	64872,
		18487	=>	64871,
		18488	=>	64871,
		18489	=>	64870,
		18490	=>	64869,
		18491	=>	64869,
		18492	=>	64868,
		18493	=>	64867,
		18494	=>	64867,
		18495	=>	64866,
		18496	=>	64866,
		18497	=>	64865,
		18498	=>	64864,
		18499	=>	64864,
		18500	=>	64863,
		18501	=>	64862,
		18502	=>	64862,
		18503	=>	64861,
		18504	=>	64860,
		18505	=>	64860,
		18506	=>	64859,
		18507	=>	64859,
		18508	=>	64858,
		18509	=>	64857,
		18510	=>	64857,
		18511	=>	64856,
		18512	=>	64855,
		18513	=>	64855,
		18514	=>	64854,
		18515	=>	64853,
		18516	=>	64853,
		18517	=>	64852,
		18518	=>	64852,
		18519	=>	64851,
		18520	=>	64850,
		18521	=>	64850,
		18522	=>	64849,
		18523	=>	64848,
		18524	=>	64848,
		18525	=>	64847,
		18526	=>	64846,
		18527	=>	64846,
		18528	=>	64845,
		18529	=>	64845,
		18530	=>	64844,
		18531	=>	64843,
		18532	=>	64843,
		18533	=>	64842,
		18534	=>	64841,
		18535	=>	64841,
		18536	=>	64840,
		18537	=>	64839,
		18538	=>	64839,
		18539	=>	64838,
		18540	=>	64837,
		18541	=>	64837,
		18542	=>	64836,
		18543	=>	64836,
		18544	=>	64835,
		18545	=>	64834,
		18546	=>	64834,
		18547	=>	64833,
		18548	=>	64832,
		18549	=>	64832,
		18550	=>	64831,
		18551	=>	64830,
		18552	=>	64830,
		18553	=>	64829,
		18554	=>	64828,
		18555	=>	64828,
		18556	=>	64827,
		18557	=>	64826,
		18558	=>	64826,
		18559	=>	64825,
		18560	=>	64825,
		18561	=>	64824,
		18562	=>	64823,
		18563	=>	64823,
		18564	=>	64822,
		18565	=>	64821,
		18566	=>	64821,
		18567	=>	64820,
		18568	=>	64819,
		18569	=>	64819,
		18570	=>	64818,
		18571	=>	64817,
		18572	=>	64817,
		18573	=>	64816,
		18574	=>	64815,
		18575	=>	64815,
		18576	=>	64814,
		18577	=>	64813,
		18578	=>	64813,
		18579	=>	64812,
		18580	=>	64811,
		18581	=>	64811,
		18582	=>	64810,
		18583	=>	64809,
		18584	=>	64809,
		18585	=>	64808,
		18586	=>	64807,
		18587	=>	64807,
		18588	=>	64806,
		18589	=>	64806,
		18590	=>	64805,
		18591	=>	64804,
		18592	=>	64804,
		18593	=>	64803,
		18594	=>	64802,
		18595	=>	64802,
		18596	=>	64801,
		18597	=>	64800,
		18598	=>	64800,
		18599	=>	64799,
		18600	=>	64798,
		18601	=>	64798,
		18602	=>	64797,
		18603	=>	64796,
		18604	=>	64796,
		18605	=>	64795,
		18606	=>	64794,
		18607	=>	64794,
		18608	=>	64793,
		18609	=>	64792,
		18610	=>	64792,
		18611	=>	64791,
		18612	=>	64790,
		18613	=>	64790,
		18614	=>	64789,
		18615	=>	64788,
		18616	=>	64788,
		18617	=>	64787,
		18618	=>	64786,
		18619	=>	64786,
		18620	=>	64785,
		18621	=>	64784,
		18622	=>	64784,
		18623	=>	64783,
		18624	=>	64782,
		18625	=>	64782,
		18626	=>	64781,
		18627	=>	64780,
		18628	=>	64780,
		18629	=>	64779,
		18630	=>	64778,
		18631	=>	64778,
		18632	=>	64777,
		18633	=>	64776,
		18634	=>	64776,
		18635	=>	64775,
		18636	=>	64774,
		18637	=>	64774,
		18638	=>	64773,
		18639	=>	64772,
		18640	=>	64772,
		18641	=>	64771,
		18642	=>	64770,
		18643	=>	64769,
		18644	=>	64769,
		18645	=>	64768,
		18646	=>	64767,
		18647	=>	64767,
		18648	=>	64766,
		18649	=>	64765,
		18650	=>	64765,
		18651	=>	64764,
		18652	=>	64763,
		18653	=>	64763,
		18654	=>	64762,
		18655	=>	64761,
		18656	=>	64761,
		18657	=>	64760,
		18658	=>	64759,
		18659	=>	64759,
		18660	=>	64758,
		18661	=>	64757,
		18662	=>	64757,
		18663	=>	64756,
		18664	=>	64755,
		18665	=>	64755,
		18666	=>	64754,
		18667	=>	64753,
		18668	=>	64753,
		18669	=>	64752,
		18670	=>	64751,
		18671	=>	64750,
		18672	=>	64750,
		18673	=>	64749,
		18674	=>	64748,
		18675	=>	64748,
		18676	=>	64747,
		18677	=>	64746,
		18678	=>	64746,
		18679	=>	64745,
		18680	=>	64744,
		18681	=>	64744,
		18682	=>	64743,
		18683	=>	64742,
		18684	=>	64742,
		18685	=>	64741,
		18686	=>	64740,
		18687	=>	64740,
		18688	=>	64739,
		18689	=>	64738,
		18690	=>	64737,
		18691	=>	64737,
		18692	=>	64736,
		18693	=>	64735,
		18694	=>	64735,
		18695	=>	64734,
		18696	=>	64733,
		18697	=>	64733,
		18698	=>	64732,
		18699	=>	64731,
		18700	=>	64731,
		18701	=>	64730,
		18702	=>	64729,
		18703	=>	64728,
		18704	=>	64728,
		18705	=>	64727,
		18706	=>	64726,
		18707	=>	64726,
		18708	=>	64725,
		18709	=>	64724,
		18710	=>	64724,
		18711	=>	64723,
		18712	=>	64722,
		18713	=>	64722,
		18714	=>	64721,
		18715	=>	64720,
		18716	=>	64719,
		18717	=>	64719,
		18718	=>	64718,
		18719	=>	64717,
		18720	=>	64717,
		18721	=>	64716,
		18722	=>	64715,
		18723	=>	64715,
		18724	=>	64714,
		18725	=>	64713,
		18726	=>	64712,
		18727	=>	64712,
		18728	=>	64711,
		18729	=>	64710,
		18730	=>	64710,
		18731	=>	64709,
		18732	=>	64708,
		18733	=>	64708,
		18734	=>	64707,
		18735	=>	64706,
		18736	=>	64705,
		18737	=>	64705,
		18738	=>	64704,
		18739	=>	64703,
		18740	=>	64703,
		18741	=>	64702,
		18742	=>	64701,
		18743	=>	64701,
		18744	=>	64700,
		18745	=>	64699,
		18746	=>	64698,
		18747	=>	64698,
		18748	=>	64697,
		18749	=>	64696,
		18750	=>	64696,
		18751	=>	64695,
		18752	=>	64694,
		18753	=>	64693,
		18754	=>	64693,
		18755	=>	64692,
		18756	=>	64691,
		18757	=>	64691,
		18758	=>	64690,
		18759	=>	64689,
		18760	=>	64688,
		18761	=>	64688,
		18762	=>	64687,
		18763	=>	64686,
		18764	=>	64686,
		18765	=>	64685,
		18766	=>	64684,
		18767	=>	64684,
		18768	=>	64683,
		18769	=>	64682,
		18770	=>	64681,
		18771	=>	64681,
		18772	=>	64680,
		18773	=>	64679,
		18774	=>	64679,
		18775	=>	64678,
		18776	=>	64677,
		18777	=>	64676,
		18778	=>	64676,
		18779	=>	64675,
		18780	=>	64674,
		18781	=>	64674,
		18782	=>	64673,
		18783	=>	64672,
		18784	=>	64671,
		18785	=>	64671,
		18786	=>	64670,
		18787	=>	64669,
		18788	=>	64669,
		18789	=>	64668,
		18790	=>	64667,
		18791	=>	64666,
		18792	=>	64666,
		18793	=>	64665,
		18794	=>	64664,
		18795	=>	64663,
		18796	=>	64663,
		18797	=>	64662,
		18798	=>	64661,
		18799	=>	64661,
		18800	=>	64660,
		18801	=>	64659,
		18802	=>	64658,
		18803	=>	64658,
		18804	=>	64657,
		18805	=>	64656,
		18806	=>	64656,
		18807	=>	64655,
		18808	=>	64654,
		18809	=>	64653,
		18810	=>	64653,
		18811	=>	64652,
		18812	=>	64651,
		18813	=>	64650,
		18814	=>	64650,
		18815	=>	64649,
		18816	=>	64648,
		18817	=>	64648,
		18818	=>	64647,
		18819	=>	64646,
		18820	=>	64645,
		18821	=>	64645,
		18822	=>	64644,
		18823	=>	64643,
		18824	=>	64642,
		18825	=>	64642,
		18826	=>	64641,
		18827	=>	64640,
		18828	=>	64640,
		18829	=>	64639,
		18830	=>	64638,
		18831	=>	64637,
		18832	=>	64637,
		18833	=>	64636,
		18834	=>	64635,
		18835	=>	64634,
		18836	=>	64634,
		18837	=>	64633,
		18838	=>	64632,
		18839	=>	64632,
		18840	=>	64631,
		18841	=>	64630,
		18842	=>	64629,
		18843	=>	64629,
		18844	=>	64628,
		18845	=>	64627,
		18846	=>	64626,
		18847	=>	64626,
		18848	=>	64625,
		18849	=>	64624,
		18850	=>	64623,
		18851	=>	64623,
		18852	=>	64622,
		18853	=>	64621,
		18854	=>	64621,
		18855	=>	64620,
		18856	=>	64619,
		18857	=>	64618,
		18858	=>	64618,
		18859	=>	64617,
		18860	=>	64616,
		18861	=>	64615,
		18862	=>	64615,
		18863	=>	64614,
		18864	=>	64613,
		18865	=>	64612,
		18866	=>	64612,
		18867	=>	64611,
		18868	=>	64610,
		18869	=>	64609,
		18870	=>	64609,
		18871	=>	64608,
		18872	=>	64607,
		18873	=>	64606,
		18874	=>	64606,
		18875	=>	64605,
		18876	=>	64604,
		18877	=>	64603,
		18878	=>	64603,
		18879	=>	64602,
		18880	=>	64601,
		18881	=>	64601,
		18882	=>	64600,
		18883	=>	64599,
		18884	=>	64598,
		18885	=>	64598,
		18886	=>	64597,
		18887	=>	64596,
		18888	=>	64595,
		18889	=>	64595,
		18890	=>	64594,
		18891	=>	64593,
		18892	=>	64592,
		18893	=>	64592,
		18894	=>	64591,
		18895	=>	64590,
		18896	=>	64589,
		18897	=>	64589,
		18898	=>	64588,
		18899	=>	64587,
		18900	=>	64586,
		18901	=>	64586,
		18902	=>	64585,
		18903	=>	64584,
		18904	=>	64583,
		18905	=>	64583,
		18906	=>	64582,
		18907	=>	64581,
		18908	=>	64580,
		18909	=>	64580,
		18910	=>	64579,
		18911	=>	64578,
		18912	=>	64577,
		18913	=>	64577,
		18914	=>	64576,
		18915	=>	64575,
		18916	=>	64574,
		18917	=>	64574,
		18918	=>	64573,
		18919	=>	64572,
		18920	=>	64571,
		18921	=>	64570,
		18922	=>	64570,
		18923	=>	64569,
		18924	=>	64568,
		18925	=>	64567,
		18926	=>	64567,
		18927	=>	64566,
		18928	=>	64565,
		18929	=>	64564,
		18930	=>	64564,
		18931	=>	64563,
		18932	=>	64562,
		18933	=>	64561,
		18934	=>	64561,
		18935	=>	64560,
		18936	=>	64559,
		18937	=>	64558,
		18938	=>	64558,
		18939	=>	64557,
		18940	=>	64556,
		18941	=>	64555,
		18942	=>	64555,
		18943	=>	64554,
		18944	=>	64553,
		18945	=>	64552,
		18946	=>	64551,
		18947	=>	64551,
		18948	=>	64550,
		18949	=>	64549,
		18950	=>	64548,
		18951	=>	64548,
		18952	=>	64547,
		18953	=>	64546,
		18954	=>	64545,
		18955	=>	64545,
		18956	=>	64544,
		18957	=>	64543,
		18958	=>	64542,
		18959	=>	64542,
		18960	=>	64541,
		18961	=>	64540,
		18962	=>	64539,
		18963	=>	64538,
		18964	=>	64538,
		18965	=>	64537,
		18966	=>	64536,
		18967	=>	64535,
		18968	=>	64535,
		18969	=>	64534,
		18970	=>	64533,
		18971	=>	64532,
		18972	=>	64532,
		18973	=>	64531,
		18974	=>	64530,
		18975	=>	64529,
		18976	=>	64528,
		18977	=>	64528,
		18978	=>	64527,
		18979	=>	64526,
		18980	=>	64525,
		18981	=>	64525,
		18982	=>	64524,
		18983	=>	64523,
		18984	=>	64522,
		18985	=>	64521,
		18986	=>	64521,
		18987	=>	64520,
		18988	=>	64519,
		18989	=>	64518,
		18990	=>	64518,
		18991	=>	64517,
		18992	=>	64516,
		18993	=>	64515,
		18994	=>	64514,
		18995	=>	64514,
		18996	=>	64513,
		18997	=>	64512,
		18998	=>	64511,
		18999	=>	64511,
		19000	=>	64510,
		19001	=>	64509,
		19002	=>	64508,
		19003	=>	64507,
		19004	=>	64507,
		19005	=>	64506,
		19006	=>	64505,
		19007	=>	64504,
		19008	=>	64504,
		19009	=>	64503,
		19010	=>	64502,
		19011	=>	64501,
		19012	=>	64500,
		19013	=>	64500,
		19014	=>	64499,
		19015	=>	64498,
		19016	=>	64497,
		19017	=>	64496,
		19018	=>	64496,
		19019	=>	64495,
		19020	=>	64494,
		19021	=>	64493,
		19022	=>	64493,
		19023	=>	64492,
		19024	=>	64491,
		19025	=>	64490,
		19026	=>	64489,
		19027	=>	64489,
		19028	=>	64488,
		19029	=>	64487,
		19030	=>	64486,
		19031	=>	64485,
		19032	=>	64485,
		19033	=>	64484,
		19034	=>	64483,
		19035	=>	64482,
		19036	=>	64482,
		19037	=>	64481,
		19038	=>	64480,
		19039	=>	64479,
		19040	=>	64478,
		19041	=>	64478,
		19042	=>	64477,
		19043	=>	64476,
		19044	=>	64475,
		19045	=>	64474,
		19046	=>	64474,
		19047	=>	64473,
		19048	=>	64472,
		19049	=>	64471,
		19050	=>	64470,
		19051	=>	64470,
		19052	=>	64469,
		19053	=>	64468,
		19054	=>	64467,
		19055	=>	64466,
		19056	=>	64466,
		19057	=>	64465,
		19058	=>	64464,
		19059	=>	64463,
		19060	=>	64462,
		19061	=>	64462,
		19062	=>	64461,
		19063	=>	64460,
		19064	=>	64459,
		19065	=>	64458,
		19066	=>	64458,
		19067	=>	64457,
		19068	=>	64456,
		19069	=>	64455,
		19070	=>	64455,
		19071	=>	64454,
		19072	=>	64453,
		19073	=>	64452,
		19074	=>	64451,
		19075	=>	64450,
		19076	=>	64450,
		19077	=>	64449,
		19078	=>	64448,
		19079	=>	64447,
		19080	=>	64446,
		19081	=>	64446,
		19082	=>	64445,
		19083	=>	64444,
		19084	=>	64443,
		19085	=>	64442,
		19086	=>	64442,
		19087	=>	64441,
		19088	=>	64440,
		19089	=>	64439,
		19090	=>	64438,
		19091	=>	64438,
		19092	=>	64437,
		19093	=>	64436,
		19094	=>	64435,
		19095	=>	64434,
		19096	=>	64434,
		19097	=>	64433,
		19098	=>	64432,
		19099	=>	64431,
		19100	=>	64430,
		19101	=>	64430,
		19102	=>	64429,
		19103	=>	64428,
		19104	=>	64427,
		19105	=>	64426,
		19106	=>	64426,
		19107	=>	64425,
		19108	=>	64424,
		19109	=>	64423,
		19110	=>	64422,
		19111	=>	64421,
		19112	=>	64421,
		19113	=>	64420,
		19114	=>	64419,
		19115	=>	64418,
		19116	=>	64417,
		19117	=>	64417,
		19118	=>	64416,
		19119	=>	64415,
		19120	=>	64414,
		19121	=>	64413,
		19122	=>	64413,
		19123	=>	64412,
		19124	=>	64411,
		19125	=>	64410,
		19126	=>	64409,
		19127	=>	64408,
		19128	=>	64408,
		19129	=>	64407,
		19130	=>	64406,
		19131	=>	64405,
		19132	=>	64404,
		19133	=>	64404,
		19134	=>	64403,
		19135	=>	64402,
		19136	=>	64401,
		19137	=>	64400,
		19138	=>	64399,
		19139	=>	64399,
		19140	=>	64398,
		19141	=>	64397,
		19142	=>	64396,
		19143	=>	64395,
		19144	=>	64394,
		19145	=>	64394,
		19146	=>	64393,
		19147	=>	64392,
		19148	=>	64391,
		19149	=>	64390,
		19150	=>	64390,
		19151	=>	64389,
		19152	=>	64388,
		19153	=>	64387,
		19154	=>	64386,
		19155	=>	64385,
		19156	=>	64385,
		19157	=>	64384,
		19158	=>	64383,
		19159	=>	64382,
		19160	=>	64381,
		19161	=>	64380,
		19162	=>	64380,
		19163	=>	64379,
		19164	=>	64378,
		19165	=>	64377,
		19166	=>	64376,
		19167	=>	64376,
		19168	=>	64375,
		19169	=>	64374,
		19170	=>	64373,
		19171	=>	64372,
		19172	=>	64371,
		19173	=>	64371,
		19174	=>	64370,
		19175	=>	64369,
		19176	=>	64368,
		19177	=>	64367,
		19178	=>	64366,
		19179	=>	64366,
		19180	=>	64365,
		19181	=>	64364,
		19182	=>	64363,
		19183	=>	64362,
		19184	=>	64361,
		19185	=>	64361,
		19186	=>	64360,
		19187	=>	64359,
		19188	=>	64358,
		19189	=>	64357,
		19190	=>	64356,
		19191	=>	64356,
		19192	=>	64355,
		19193	=>	64354,
		19194	=>	64353,
		19195	=>	64352,
		19196	=>	64351,
		19197	=>	64351,
		19198	=>	64350,
		19199	=>	64349,
		19200	=>	64348,
		19201	=>	64347,
		19202	=>	64346,
		19203	=>	64346,
		19204	=>	64345,
		19205	=>	64344,
		19206	=>	64343,
		19207	=>	64342,
		19208	=>	64341,
		19209	=>	64340,
		19210	=>	64340,
		19211	=>	64339,
		19212	=>	64338,
		19213	=>	64337,
		19214	=>	64336,
		19215	=>	64335,
		19216	=>	64335,
		19217	=>	64334,
		19218	=>	64333,
		19219	=>	64332,
		19220	=>	64331,
		19221	=>	64330,
		19222	=>	64330,
		19223	=>	64329,
		19224	=>	64328,
		19225	=>	64327,
		19226	=>	64326,
		19227	=>	64325,
		19228	=>	64324,
		19229	=>	64324,
		19230	=>	64323,
		19231	=>	64322,
		19232	=>	64321,
		19233	=>	64320,
		19234	=>	64319,
		19235	=>	64319,
		19236	=>	64318,
		19237	=>	64317,
		19238	=>	64316,
		19239	=>	64315,
		19240	=>	64314,
		19241	=>	64313,
		19242	=>	64313,
		19243	=>	64312,
		19244	=>	64311,
		19245	=>	64310,
		19246	=>	64309,
		19247	=>	64308,
		19248	=>	64307,
		19249	=>	64307,
		19250	=>	64306,
		19251	=>	64305,
		19252	=>	64304,
		19253	=>	64303,
		19254	=>	64302,
		19255	=>	64302,
		19256	=>	64301,
		19257	=>	64300,
		19258	=>	64299,
		19259	=>	64298,
		19260	=>	64297,
		19261	=>	64296,
		19262	=>	64296,
		19263	=>	64295,
		19264	=>	64294,
		19265	=>	64293,
		19266	=>	64292,
		19267	=>	64291,
		19268	=>	64290,
		19269	=>	64290,
		19270	=>	64289,
		19271	=>	64288,
		19272	=>	64287,
		19273	=>	64286,
		19274	=>	64285,
		19275	=>	64284,
		19276	=>	64284,
		19277	=>	64283,
		19278	=>	64282,
		19279	=>	64281,
		19280	=>	64280,
		19281	=>	64279,
		19282	=>	64278,
		19283	=>	64277,
		19284	=>	64277,
		19285	=>	64276,
		19286	=>	64275,
		19287	=>	64274,
		19288	=>	64273,
		19289	=>	64272,
		19290	=>	64271,
		19291	=>	64271,
		19292	=>	64270,
		19293	=>	64269,
		19294	=>	64268,
		19295	=>	64267,
		19296	=>	64266,
		19297	=>	64265,
		19298	=>	64265,
		19299	=>	64264,
		19300	=>	64263,
		19301	=>	64262,
		19302	=>	64261,
		19303	=>	64260,
		19304	=>	64259,
		19305	=>	64258,
		19306	=>	64258,
		19307	=>	64257,
		19308	=>	64256,
		19309	=>	64255,
		19310	=>	64254,
		19311	=>	64253,
		19312	=>	64252,
		19313	=>	64251,
		19314	=>	64251,
		19315	=>	64250,
		19316	=>	64249,
		19317	=>	64248,
		19318	=>	64247,
		19319	=>	64246,
		19320	=>	64245,
		19321	=>	64245,
		19322	=>	64244,
		19323	=>	64243,
		19324	=>	64242,
		19325	=>	64241,
		19326	=>	64240,
		19327	=>	64239,
		19328	=>	64238,
		19329	=>	64238,
		19330	=>	64237,
		19331	=>	64236,
		19332	=>	64235,
		19333	=>	64234,
		19334	=>	64233,
		19335	=>	64232,
		19336	=>	64231,
		19337	=>	64231,
		19338	=>	64230,
		19339	=>	64229,
		19340	=>	64228,
		19341	=>	64227,
		19342	=>	64226,
		19343	=>	64225,
		19344	=>	64224,
		19345	=>	64223,
		19346	=>	64223,
		19347	=>	64222,
		19348	=>	64221,
		19349	=>	64220,
		19350	=>	64219,
		19351	=>	64218,
		19352	=>	64217,
		19353	=>	64216,
		19354	=>	64216,
		19355	=>	64215,
		19356	=>	64214,
		19357	=>	64213,
		19358	=>	64212,
		19359	=>	64211,
		19360	=>	64210,
		19361	=>	64209,
		19362	=>	64208,
		19363	=>	64208,
		19364	=>	64207,
		19365	=>	64206,
		19366	=>	64205,
		19367	=>	64204,
		19368	=>	64203,
		19369	=>	64202,
		19370	=>	64201,
		19371	=>	64201,
		19372	=>	64200,
		19373	=>	64199,
		19374	=>	64198,
		19375	=>	64197,
		19376	=>	64196,
		19377	=>	64195,
		19378	=>	64194,
		19379	=>	64193,
		19380	=>	64193,
		19381	=>	64192,
		19382	=>	64191,
		19383	=>	64190,
		19384	=>	64189,
		19385	=>	64188,
		19386	=>	64187,
		19387	=>	64186,
		19388	=>	64185,
		19389	=>	64184,
		19390	=>	64184,
		19391	=>	64183,
		19392	=>	64182,
		19393	=>	64181,
		19394	=>	64180,
		19395	=>	64179,
		19396	=>	64178,
		19397	=>	64177,
		19398	=>	64176,
		19399	=>	64176,
		19400	=>	64175,
		19401	=>	64174,
		19402	=>	64173,
		19403	=>	64172,
		19404	=>	64171,
		19405	=>	64170,
		19406	=>	64169,
		19407	=>	64168,
		19408	=>	64167,
		19409	=>	64167,
		19410	=>	64166,
		19411	=>	64165,
		19412	=>	64164,
		19413	=>	64163,
		19414	=>	64162,
		19415	=>	64161,
		19416	=>	64160,
		19417	=>	64159,
		19418	=>	64158,
		19419	=>	64158,
		19420	=>	64157,
		19421	=>	64156,
		19422	=>	64155,
		19423	=>	64154,
		19424	=>	64153,
		19425	=>	64152,
		19426	=>	64151,
		19427	=>	64150,
		19428	=>	64149,
		19429	=>	64149,
		19430	=>	64148,
		19431	=>	64147,
		19432	=>	64146,
		19433	=>	64145,
		19434	=>	64144,
		19435	=>	64143,
		19436	=>	64142,
		19437	=>	64141,
		19438	=>	64140,
		19439	=>	64140,
		19440	=>	64139,
		19441	=>	64138,
		19442	=>	64137,
		19443	=>	64136,
		19444	=>	64135,
		19445	=>	64134,
		19446	=>	64133,
		19447	=>	64132,
		19448	=>	64131,
		19449	=>	64130,
		19450	=>	64130,
		19451	=>	64129,
		19452	=>	64128,
		19453	=>	64127,
		19454	=>	64126,
		19455	=>	64125,
		19456	=>	64124,
		19457	=>	64123,
		19458	=>	64122,
		19459	=>	64121,
		19460	=>	64120,
		19461	=>	64119,
		19462	=>	64119,
		19463	=>	64118,
		19464	=>	64117,
		19465	=>	64116,
		19466	=>	64115,
		19467	=>	64114,
		19468	=>	64113,
		19469	=>	64112,
		19470	=>	64111,
		19471	=>	64110,
		19472	=>	64109,
		19473	=>	64108,
		19474	=>	64108,
		19475	=>	64107,
		19476	=>	64106,
		19477	=>	64105,
		19478	=>	64104,
		19479	=>	64103,
		19480	=>	64102,
		19481	=>	64101,
		19482	=>	64100,
		19483	=>	64099,
		19484	=>	64098,
		19485	=>	64097,
		19486	=>	64097,
		19487	=>	64096,
		19488	=>	64095,
		19489	=>	64094,
		19490	=>	64093,
		19491	=>	64092,
		19492	=>	64091,
		19493	=>	64090,
		19494	=>	64089,
		19495	=>	64088,
		19496	=>	64087,
		19497	=>	64086,
		19498	=>	64085,
		19499	=>	64085,
		19500	=>	64084,
		19501	=>	64083,
		19502	=>	64082,
		19503	=>	64081,
		19504	=>	64080,
		19505	=>	64079,
		19506	=>	64078,
		19507	=>	64077,
		19508	=>	64076,
		19509	=>	64075,
		19510	=>	64074,
		19511	=>	64073,
		19512	=>	64073,
		19513	=>	64072,
		19514	=>	64071,
		19515	=>	64070,
		19516	=>	64069,
		19517	=>	64068,
		19518	=>	64067,
		19519	=>	64066,
		19520	=>	64065,
		19521	=>	64064,
		19522	=>	64063,
		19523	=>	64062,
		19524	=>	64061,
		19525	=>	64060,
		19526	=>	64060,
		19527	=>	64059,
		19528	=>	64058,
		19529	=>	64057,
		19530	=>	64056,
		19531	=>	64055,
		19532	=>	64054,
		19533	=>	64053,
		19534	=>	64052,
		19535	=>	64051,
		19536	=>	64050,
		19537	=>	64049,
		19538	=>	64048,
		19539	=>	64047,
		19540	=>	64046,
		19541	=>	64045,
		19542	=>	64045,
		19543	=>	64044,
		19544	=>	64043,
		19545	=>	64042,
		19546	=>	64041,
		19547	=>	64040,
		19548	=>	64039,
		19549	=>	64038,
		19550	=>	64037,
		19551	=>	64036,
		19552	=>	64035,
		19553	=>	64034,
		19554	=>	64033,
		19555	=>	64032,
		19556	=>	64031,
		19557	=>	64030,
		19558	=>	64030,
		19559	=>	64029,
		19560	=>	64028,
		19561	=>	64027,
		19562	=>	64026,
		19563	=>	64025,
		19564	=>	64024,
		19565	=>	64023,
		19566	=>	64022,
		19567	=>	64021,
		19568	=>	64020,
		19569	=>	64019,
		19570	=>	64018,
		19571	=>	64017,
		19572	=>	64016,
		19573	=>	64015,
		19574	=>	64014,
		19575	=>	64013,
		19576	=>	64013,
		19577	=>	64012,
		19578	=>	64011,
		19579	=>	64010,
		19580	=>	64009,
		19581	=>	64008,
		19582	=>	64007,
		19583	=>	64006,
		19584	=>	64005,
		19585	=>	64004,
		19586	=>	64003,
		19587	=>	64002,
		19588	=>	64001,
		19589	=>	64000,
		19590	=>	63999,
		19591	=>	63998,
		19592	=>	63997,
		19593	=>	63996,
		19594	=>	63995,
		19595	=>	63995,
		19596	=>	63994,
		19597	=>	63993,
		19598	=>	63992,
		19599	=>	63991,
		19600	=>	63990,
		19601	=>	63989,
		19602	=>	63988,
		19603	=>	63987,
		19604	=>	63986,
		19605	=>	63985,
		19606	=>	63984,
		19607	=>	63983,
		19608	=>	63982,
		19609	=>	63981,
		19610	=>	63980,
		19611	=>	63979,
		19612	=>	63978,
		19613	=>	63977,
		19614	=>	63976,
		19615	=>	63975,
		19616	=>	63974,
		19617	=>	63973,
		19618	=>	63973,
		19619	=>	63972,
		19620	=>	63971,
		19621	=>	63970,
		19622	=>	63969,
		19623	=>	63968,
		19624	=>	63967,
		19625	=>	63966,
		19626	=>	63965,
		19627	=>	63964,
		19628	=>	63963,
		19629	=>	63962,
		19630	=>	63961,
		19631	=>	63960,
		19632	=>	63959,
		19633	=>	63958,
		19634	=>	63957,
		19635	=>	63956,
		19636	=>	63955,
		19637	=>	63954,
		19638	=>	63953,
		19639	=>	63952,
		19640	=>	63951,
		19641	=>	63950,
		19642	=>	63949,
		19643	=>	63948,
		19644	=>	63948,
		19645	=>	63947,
		19646	=>	63946,
		19647	=>	63945,
		19648	=>	63944,
		19649	=>	63943,
		19650	=>	63942,
		19651	=>	63941,
		19652	=>	63940,
		19653	=>	63939,
		19654	=>	63938,
		19655	=>	63937,
		19656	=>	63936,
		19657	=>	63935,
		19658	=>	63934,
		19659	=>	63933,
		19660	=>	63932,
		19661	=>	63931,
		19662	=>	63930,
		19663	=>	63929,
		19664	=>	63928,
		19665	=>	63927,
		19666	=>	63926,
		19667	=>	63925,
		19668	=>	63924,
		19669	=>	63923,
		19670	=>	63922,
		19671	=>	63921,
		19672	=>	63920,
		19673	=>	63919,
		19674	=>	63918,
		19675	=>	63917,
		19676	=>	63916,
		19677	=>	63915,
		19678	=>	63915,
		19679	=>	63914,
		19680	=>	63913,
		19681	=>	63912,
		19682	=>	63911,
		19683	=>	63910,
		19684	=>	63909,
		19685	=>	63908,
		19686	=>	63907,
		19687	=>	63906,
		19688	=>	63905,
		19689	=>	63904,
		19690	=>	63903,
		19691	=>	63902,
		19692	=>	63901,
		19693	=>	63900,
		19694	=>	63899,
		19695	=>	63898,
		19696	=>	63897,
		19697	=>	63896,
		19698	=>	63895,
		19699	=>	63894,
		19700	=>	63893,
		19701	=>	63892,
		19702	=>	63891,
		19703	=>	63890,
		19704	=>	63889,
		19705	=>	63888,
		19706	=>	63887,
		19707	=>	63886,
		19708	=>	63885,
		19709	=>	63884,
		19710	=>	63883,
		19711	=>	63882,
		19712	=>	63881,
		19713	=>	63880,
		19714	=>	63879,
		19715	=>	63878,
		19716	=>	63877,
		19717	=>	63876,
		19718	=>	63875,
		19719	=>	63874,
		19720	=>	63873,
		19721	=>	63872,
		19722	=>	63871,
		19723	=>	63870,
		19724	=>	63869,
		19725	=>	63868,
		19726	=>	63867,
		19727	=>	63866,
		19728	=>	63865,
		19729	=>	63864,
		19730	=>	63863,
		19731	=>	63862,
		19732	=>	63861,
		19733	=>	63860,
		19734	=>	63859,
		19735	=>	63858,
		19736	=>	63857,
		19737	=>	63856,
		19738	=>	63855,
		19739	=>	63854,
		19740	=>	63853,
		19741	=>	63852,
		19742	=>	63851,
		19743	=>	63850,
		19744	=>	63849,
		19745	=>	63848,
		19746	=>	63847,
		19747	=>	63846,
		19748	=>	63846,
		19749	=>	63845,
		19750	=>	63844,
		19751	=>	63843,
		19752	=>	63842,
		19753	=>	63841,
		19754	=>	63840,
		19755	=>	63839,
		19756	=>	63838,
		19757	=>	63837,
		19758	=>	63836,
		19759	=>	63835,
		19760	=>	63834,
		19761	=>	63833,
		19762	=>	63832,
		19763	=>	63831,
		19764	=>	63830,
		19765	=>	63829,
		19766	=>	63828,
		19767	=>	63827,
		19768	=>	63826,
		19769	=>	63825,
		19770	=>	63824,
		19771	=>	63823,
		19772	=>	63822,
		19773	=>	63821,
		19774	=>	63820,
		19775	=>	63819,
		19776	=>	63818,
		19777	=>	63817,
		19778	=>	63816,
		19779	=>	63814,
		19780	=>	63813,
		19781	=>	63812,
		19782	=>	63811,
		19783	=>	63810,
		19784	=>	63809,
		19785	=>	63808,
		19786	=>	63807,
		19787	=>	63806,
		19788	=>	63805,
		19789	=>	63804,
		19790	=>	63803,
		19791	=>	63802,
		19792	=>	63801,
		19793	=>	63800,
		19794	=>	63799,
		19795	=>	63798,
		19796	=>	63797,
		19797	=>	63796,
		19798	=>	63795,
		19799	=>	63794,
		19800	=>	63793,
		19801	=>	63792,
		19802	=>	63791,
		19803	=>	63790,
		19804	=>	63789,
		19805	=>	63788,
		19806	=>	63787,
		19807	=>	63786,
		19808	=>	63785,
		19809	=>	63784,
		19810	=>	63783,
		19811	=>	63782,
		19812	=>	63781,
		19813	=>	63780,
		19814	=>	63779,
		19815	=>	63778,
		19816	=>	63777,
		19817	=>	63776,
		19818	=>	63775,
		19819	=>	63774,
		19820	=>	63773,
		19821	=>	63772,
		19822	=>	63771,
		19823	=>	63770,
		19824	=>	63769,
		19825	=>	63768,
		19826	=>	63767,
		19827	=>	63766,
		19828	=>	63765,
		19829	=>	63764,
		19830	=>	63763,
		19831	=>	63762,
		19832	=>	63761,
		19833	=>	63760,
		19834	=>	63759,
		19835	=>	63758,
		19836	=>	63757,
		19837	=>	63756,
		19838	=>	63755,
		19839	=>	63754,
		19840	=>	63753,
		19841	=>	63752,
		19842	=>	63751,
		19843	=>	63750,
		19844	=>	63749,
		19845	=>	63748,
		19846	=>	63747,
		19847	=>	63746,
		19848	=>	63745,
		19849	=>	63743,
		19850	=>	63742,
		19851	=>	63741,
		19852	=>	63740,
		19853	=>	63739,
		19854	=>	63738,
		19855	=>	63737,
		19856	=>	63736,
		19857	=>	63735,
		19858	=>	63734,
		19859	=>	63733,
		19860	=>	63732,
		19861	=>	63731,
		19862	=>	63730,
		19863	=>	63729,
		19864	=>	63728,
		19865	=>	63727,
		19866	=>	63726,
		19867	=>	63725,
		19868	=>	63724,
		19869	=>	63723,
		19870	=>	63722,
		19871	=>	63721,
		19872	=>	63720,
		19873	=>	63719,
		19874	=>	63718,
		19875	=>	63717,
		19876	=>	63716,
		19877	=>	63715,
		19878	=>	63714,
		19879	=>	63713,
		19880	=>	63712,
		19881	=>	63711,
		19882	=>	63710,
		19883	=>	63708,
		19884	=>	63707,
		19885	=>	63706,
		19886	=>	63705,
		19887	=>	63704,
		19888	=>	63703,
		19889	=>	63702,
		19890	=>	63701,
		19891	=>	63700,
		19892	=>	63699,
		19893	=>	63698,
		19894	=>	63697,
		19895	=>	63696,
		19896	=>	63695,
		19897	=>	63694,
		19898	=>	63693,
		19899	=>	63692,
		19900	=>	63691,
		19901	=>	63690,
		19902	=>	63689,
		19903	=>	63688,
		19904	=>	63687,
		19905	=>	63686,
		19906	=>	63685,
		19907	=>	63684,
		19908	=>	63683,
		19909	=>	63681,
		19910	=>	63680,
		19911	=>	63679,
		19912	=>	63678,
		19913	=>	63677,
		19914	=>	63676,
		19915	=>	63675,
		19916	=>	63674,
		19917	=>	63673,
		19918	=>	63672,
		19919	=>	63671,
		19920	=>	63670,
		19921	=>	63669,
		19922	=>	63668,
		19923	=>	63667,
		19924	=>	63666,
		19925	=>	63665,
		19926	=>	63664,
		19927	=>	63663,
		19928	=>	63662,
		19929	=>	63661,
		19930	=>	63660,
		19931	=>	63659,
		19932	=>	63657,
		19933	=>	63656,
		19934	=>	63655,
		19935	=>	63654,
		19936	=>	63653,
		19937	=>	63652,
		19938	=>	63651,
		19939	=>	63650,
		19940	=>	63649,
		19941	=>	63648,
		19942	=>	63647,
		19943	=>	63646,
		19944	=>	63645,
		19945	=>	63644,
		19946	=>	63643,
		19947	=>	63642,
		19948	=>	63641,
		19949	=>	63640,
		19950	=>	63639,
		19951	=>	63637,
		19952	=>	63636,
		19953	=>	63635,
		19954	=>	63634,
		19955	=>	63633,
		19956	=>	63632,
		19957	=>	63631,
		19958	=>	63630,
		19959	=>	63629,
		19960	=>	63628,
		19961	=>	63627,
		19962	=>	63626,
		19963	=>	63625,
		19964	=>	63624,
		19965	=>	63623,
		19966	=>	63622,
		19967	=>	63621,
		19968	=>	63620,
		19969	=>	63618,
		19970	=>	63617,
		19971	=>	63616,
		19972	=>	63615,
		19973	=>	63614,
		19974	=>	63613,
		19975	=>	63612,
		19976	=>	63611,
		19977	=>	63610,
		19978	=>	63609,
		19979	=>	63608,
		19980	=>	63607,
		19981	=>	63606,
		19982	=>	63605,
		19983	=>	63604,
		19984	=>	63603,
		19985	=>	63602,
		19986	=>	63600,
		19987	=>	63599,
		19988	=>	63598,
		19989	=>	63597,
		19990	=>	63596,
		19991	=>	63595,
		19992	=>	63594,
		19993	=>	63593,
		19994	=>	63592,
		19995	=>	63591,
		19996	=>	63590,
		19997	=>	63589,
		19998	=>	63588,
		19999	=>	63587,
		20000	=>	63586,
		20001	=>	63584,
		20002	=>	63583,
		20003	=>	63582,
		20004	=>	63581,
		20005	=>	63580,
		20006	=>	63579,
		20007	=>	63578,
		20008	=>	63577,
		20009	=>	63576,
		20010	=>	63575,
		20011	=>	63574,
		20012	=>	63573,
		20013	=>	63572,
		20014	=>	63571,
		20015	=>	63569,
		20016	=>	63568,
		20017	=>	63567,
		20018	=>	63566,
		20019	=>	63565,
		20020	=>	63564,
		20021	=>	63563,
		20022	=>	63562,
		20023	=>	63561,
		20024	=>	63560,
		20025	=>	63559,
		20026	=>	63558,
		20027	=>	63557,
		20028	=>	63556,
		20029	=>	63554,
		20030	=>	63553,
		20031	=>	63552,
		20032	=>	63551,
		20033	=>	63550,
		20034	=>	63549,
		20035	=>	63548,
		20036	=>	63547,
		20037	=>	63546,
		20038	=>	63545,
		20039	=>	63544,
		20040	=>	63543,
		20041	=>	63542,
		20042	=>	63540,
		20043	=>	63539,
		20044	=>	63538,
		20045	=>	63537,
		20046	=>	63536,
		20047	=>	63535,
		20048	=>	63534,
		20049	=>	63533,
		20050	=>	63532,
		20051	=>	63531,
		20052	=>	63530,
		20053	=>	63529,
		20054	=>	63527,
		20055	=>	63526,
		20056	=>	63525,
		20057	=>	63524,
		20058	=>	63523,
		20059	=>	63522,
		20060	=>	63521,
		20061	=>	63520,
		20062	=>	63519,
		20063	=>	63518,
		20064	=>	63517,
		20065	=>	63516,
		20066	=>	63514,
		20067	=>	63513,
		20068	=>	63512,
		20069	=>	63511,
		20070	=>	63510,
		20071	=>	63509,
		20072	=>	63508,
		20073	=>	63507,
		20074	=>	63506,
		20075	=>	63505,
		20076	=>	63504,
		20077	=>	63503,
		20078	=>	63501,
		20079	=>	63500,
		20080	=>	63499,
		20081	=>	63498,
		20082	=>	63497,
		20083	=>	63496,
		20084	=>	63495,
		20085	=>	63494,
		20086	=>	63493,
		20087	=>	63492,
		20088	=>	63491,
		20089	=>	63489,
		20090	=>	63488,
		20091	=>	63487,
		20092	=>	63486,
		20093	=>	63485,
		20094	=>	63484,
		20095	=>	63483,
		20096	=>	63482,
		20097	=>	63481,
		20098	=>	63480,
		20099	=>	63478,
		20100	=>	63477,
		20101	=>	63476,
		20102	=>	63475,
		20103	=>	63474,
		20104	=>	63473,
		20105	=>	63472,
		20106	=>	63471,
		20107	=>	63470,
		20108	=>	63469,
		20109	=>	63468,
		20110	=>	63466,
		20111	=>	63465,
		20112	=>	63464,
		20113	=>	63463,
		20114	=>	63462,
		20115	=>	63461,
		20116	=>	63460,
		20117	=>	63459,
		20118	=>	63458,
		20119	=>	63457,
		20120	=>	63455,
		20121	=>	63454,
		20122	=>	63453,
		20123	=>	63452,
		20124	=>	63451,
		20125	=>	63450,
		20126	=>	63449,
		20127	=>	63448,
		20128	=>	63447,
		20129	=>	63445,
		20130	=>	63444,
		20131	=>	63443,
		20132	=>	63442,
		20133	=>	63441,
		20134	=>	63440,
		20135	=>	63439,
		20136	=>	63438,
		20137	=>	63437,
		20138	=>	63436,
		20139	=>	63434,
		20140	=>	63433,
		20141	=>	63432,
		20142	=>	63431,
		20143	=>	63430,
		20144	=>	63429,
		20145	=>	63428,
		20146	=>	63427,
		20147	=>	63426,
		20148	=>	63424,
		20149	=>	63423,
		20150	=>	63422,
		20151	=>	63421,
		20152	=>	63420,
		20153	=>	63419,
		20154	=>	63418,
		20155	=>	63417,
		20156	=>	63416,
		20157	=>	63414,
		20158	=>	63413,
		20159	=>	63412,
		20160	=>	63411,
		20161	=>	63410,
		20162	=>	63409,
		20163	=>	63408,
		20164	=>	63407,
		20165	=>	63406,
		20166	=>	63404,
		20167	=>	63403,
		20168	=>	63402,
		20169	=>	63401,
		20170	=>	63400,
		20171	=>	63399,
		20172	=>	63398,
		20173	=>	63397,
		20174	=>	63396,
		20175	=>	63394,
		20176	=>	63393,
		20177	=>	63392,
		20178	=>	63391,
		20179	=>	63390,
		20180	=>	63389,
		20181	=>	63388,
		20182	=>	63387,
		20183	=>	63385,
		20184	=>	63384,
		20185	=>	63383,
		20186	=>	63382,
		20187	=>	63381,
		20188	=>	63380,
		20189	=>	63379,
		20190	=>	63378,
		20191	=>	63376,
		20192	=>	63375,
		20193	=>	63374,
		20194	=>	63373,
		20195	=>	63372,
		20196	=>	63371,
		20197	=>	63370,
		20198	=>	63369,
		20199	=>	63368,
		20200	=>	63366,
		20201	=>	63365,
		20202	=>	63364,
		20203	=>	63363,
		20204	=>	63362,
		20205	=>	63361,
		20206	=>	63360,
		20207	=>	63359,
		20208	=>	63357,
		20209	=>	63356,
		20210	=>	63355,
		20211	=>	63354,
		20212	=>	63353,
		20213	=>	63352,
		20214	=>	63351,
		20215	=>	63350,
		20216	=>	63348,
		20217	=>	63347,
		20218	=>	63346,
		20219	=>	63345,
		20220	=>	63344,
		20221	=>	63343,
		20222	=>	63342,
		20223	=>	63340,
		20224	=>	63339,
		20225	=>	63338,
		20226	=>	63337,
		20227	=>	63336,
		20228	=>	63335,
		20229	=>	63334,
		20230	=>	63333,
		20231	=>	63331,
		20232	=>	63330,
		20233	=>	63329,
		20234	=>	63328,
		20235	=>	63327,
		20236	=>	63326,
		20237	=>	63325,
		20238	=>	63323,
		20239	=>	63322,
		20240	=>	63321,
		20241	=>	63320,
		20242	=>	63319,
		20243	=>	63318,
		20244	=>	63317,
		20245	=>	63316,
		20246	=>	63314,
		20247	=>	63313,
		20248	=>	63312,
		20249	=>	63311,
		20250	=>	63310,
		20251	=>	63309,
		20252	=>	63308,
		20253	=>	63306,
		20254	=>	63305,
		20255	=>	63304,
		20256	=>	63303,
		20257	=>	63302,
		20258	=>	63301,
		20259	=>	63300,
		20260	=>	63298,
		20261	=>	63297,
		20262	=>	63296,
		20263	=>	63295,
		20264	=>	63294,
		20265	=>	63293,
		20266	=>	63292,
		20267	=>	63290,
		20268	=>	63289,
		20269	=>	63288,
		20270	=>	63287,
		20271	=>	63286,
		20272	=>	63285,
		20273	=>	63284,
		20274	=>	63282,
		20275	=>	63281,
		20276	=>	63280,
		20277	=>	63279,
		20278	=>	63278,
		20279	=>	63277,
		20280	=>	63276,
		20281	=>	63274,
		20282	=>	63273,
		20283	=>	63272,
		20284	=>	63271,
		20285	=>	63270,
		20286	=>	63269,
		20287	=>	63268,
		20288	=>	63266,
		20289	=>	63265,
		20290	=>	63264,
		20291	=>	63263,
		20292	=>	63262,
		20293	=>	63261,
		20294	=>	63260,
		20295	=>	63258,
		20296	=>	63257,
		20297	=>	63256,
		20298	=>	63255,
		20299	=>	63254,
		20300	=>	63253,
		20301	=>	63251,
		20302	=>	63250,
		20303	=>	63249,
		20304	=>	63248,
		20305	=>	63247,
		20306	=>	63246,
		20307	=>	63245,
		20308	=>	63243,
		20309	=>	63242,
		20310	=>	63241,
		20311	=>	63240,
		20312	=>	63239,
		20313	=>	63238,
		20314	=>	63236,
		20315	=>	63235,
		20316	=>	63234,
		20317	=>	63233,
		20318	=>	63232,
		20319	=>	63231,
		20320	=>	63230,
		20321	=>	63228,
		20322	=>	63227,
		20323	=>	63226,
		20324	=>	63225,
		20325	=>	63224,
		20326	=>	63223,
		20327	=>	63221,
		20328	=>	63220,
		20329	=>	63219,
		20330	=>	63218,
		20331	=>	63217,
		20332	=>	63216,
		20333	=>	63214,
		20334	=>	63213,
		20335	=>	63212,
		20336	=>	63211,
		20337	=>	63210,
		20338	=>	63209,
		20339	=>	63207,
		20340	=>	63206,
		20341	=>	63205,
		20342	=>	63204,
		20343	=>	63203,
		20344	=>	63202,
		20345	=>	63200,
		20346	=>	63199,
		20347	=>	63198,
		20348	=>	63197,
		20349	=>	63196,
		20350	=>	63195,
		20351	=>	63193,
		20352	=>	63192,
		20353	=>	63191,
		20354	=>	63190,
		20355	=>	63189,
		20356	=>	63188,
		20357	=>	63186,
		20358	=>	63185,
		20359	=>	63184,
		20360	=>	63183,
		20361	=>	63182,
		20362	=>	63181,
		20363	=>	63179,
		20364	=>	63178,
		20365	=>	63177,
		20366	=>	63176,
		20367	=>	63175,
		20368	=>	63174,
		20369	=>	63172,
		20370	=>	63171,
		20371	=>	63170,
		20372	=>	63169,
		20373	=>	63168,
		20374	=>	63167,
		20375	=>	63165,
		20376	=>	63164,
		20377	=>	63163,
		20378	=>	63162,
		20379	=>	63161,
		20380	=>	63160,
		20381	=>	63158,
		20382	=>	63157,
		20383	=>	63156,
		20384	=>	63155,
		20385	=>	63154,
		20386	=>	63153,
		20387	=>	63151,
		20388	=>	63150,
		20389	=>	63149,
		20390	=>	63148,
		20391	=>	63147,
		20392	=>	63145,
		20393	=>	63144,
		20394	=>	63143,
		20395	=>	63142,
		20396	=>	63141,
		20397	=>	63140,
		20398	=>	63138,
		20399	=>	63137,
		20400	=>	63136,
		20401	=>	63135,
		20402	=>	63134,
		20403	=>	63132,
		20404	=>	63131,
		20405	=>	63130,
		20406	=>	63129,
		20407	=>	63128,
		20408	=>	63127,
		20409	=>	63125,
		20410	=>	63124,
		20411	=>	63123,
		20412	=>	63122,
		20413	=>	63121,
		20414	=>	63119,
		20415	=>	63118,
		20416	=>	63117,
		20417	=>	63116,
		20418	=>	63115,
		20419	=>	63114,
		20420	=>	63112,
		20421	=>	63111,
		20422	=>	63110,
		20423	=>	63109,
		20424	=>	63108,
		20425	=>	63106,
		20426	=>	63105,
		20427	=>	63104,
		20428	=>	63103,
		20429	=>	63102,
		20430	=>	63100,
		20431	=>	63099,
		20432	=>	63098,
		20433	=>	63097,
		20434	=>	63096,
		20435	=>	63095,
		20436	=>	63093,
		20437	=>	63092,
		20438	=>	63091,
		20439	=>	63090,
		20440	=>	63089,
		20441	=>	63087,
		20442	=>	63086,
		20443	=>	63085,
		20444	=>	63084,
		20445	=>	63083,
		20446	=>	63081,
		20447	=>	63080,
		20448	=>	63079,
		20449	=>	63078,
		20450	=>	63077,
		20451	=>	63075,
		20452	=>	63074,
		20453	=>	63073,
		20454	=>	63072,
		20455	=>	63071,
		20456	=>	63069,
		20457	=>	63068,
		20458	=>	63067,
		20459	=>	63066,
		20460	=>	63065,
		20461	=>	63064,
		20462	=>	63062,
		20463	=>	63061,
		20464	=>	63060,
		20465	=>	63059,
		20466	=>	63058,
		20467	=>	63056,
		20468	=>	63055,
		20469	=>	63054,
		20470	=>	63053,
		20471	=>	63052,
		20472	=>	63050,
		20473	=>	63049,
		20474	=>	63048,
		20475	=>	63047,
		20476	=>	63046,
		20477	=>	63044,
		20478	=>	63043,
		20479	=>	63042,
		20480	=>	63041,
		20481	=>	63040,
		20482	=>	63038,
		20483	=>	63037,
		20484	=>	63036,
		20485	=>	63035,
		20486	=>	63034,
		20487	=>	63032,
		20488	=>	63031,
		20489	=>	63030,
		20490	=>	63029,
		20491	=>	63027,
		20492	=>	63026,
		20493	=>	63025,
		20494	=>	63024,
		20495	=>	63023,
		20496	=>	63021,
		20497	=>	63020,
		20498	=>	63019,
		20499	=>	63018,
		20500	=>	63017,
		20501	=>	63015,
		20502	=>	63014,
		20503	=>	63013,
		20504	=>	63012,
		20505	=>	63011,
		20506	=>	63009,
		20507	=>	63008,
		20508	=>	63007,
		20509	=>	63006,
		20510	=>	63005,
		20511	=>	63003,
		20512	=>	63002,
		20513	=>	63001,
		20514	=>	63000,
		20515	=>	62998,
		20516	=>	62997,
		20517	=>	62996,
		20518	=>	62995,
		20519	=>	62994,
		20520	=>	62992,
		20521	=>	62991,
		20522	=>	62990,
		20523	=>	62989,
		20524	=>	62988,
		20525	=>	62986,
		20526	=>	62985,
		20527	=>	62984,
		20528	=>	62983,
		20529	=>	62981,
		20530	=>	62980,
		20531	=>	62979,
		20532	=>	62978,
		20533	=>	62977,
		20534	=>	62975,
		20535	=>	62974,
		20536	=>	62973,
		20537	=>	62972,
		20538	=>	62971,
		20539	=>	62969,
		20540	=>	62968,
		20541	=>	62967,
		20542	=>	62966,
		20543	=>	62964,
		20544	=>	62963,
		20545	=>	62962,
		20546	=>	62961,
		20547	=>	62960,
		20548	=>	62958,
		20549	=>	62957,
		20550	=>	62956,
		20551	=>	62955,
		20552	=>	62953,
		20553	=>	62952,
		20554	=>	62951,
		20555	=>	62950,
		20556	=>	62949,
		20557	=>	62947,
		20558	=>	62946,
		20559	=>	62945,
		20560	=>	62944,
		20561	=>	62942,
		20562	=>	62941,
		20563	=>	62940,
		20564	=>	62939,
		20565	=>	62938,
		20566	=>	62936,
		20567	=>	62935,
		20568	=>	62934,
		20569	=>	62933,
		20570	=>	62931,
		20571	=>	62930,
		20572	=>	62929,
		20573	=>	62928,
		20574	=>	62926,
		20575	=>	62925,
		20576	=>	62924,
		20577	=>	62923,
		20578	=>	62922,
		20579	=>	62920,
		20580	=>	62919,
		20581	=>	62918,
		20582	=>	62917,
		20583	=>	62915,
		20584	=>	62914,
		20585	=>	62913,
		20586	=>	62912,
		20587	=>	62910,
		20588	=>	62909,
		20589	=>	62908,
		20590	=>	62907,
		20591	=>	62906,
		20592	=>	62904,
		20593	=>	62903,
		20594	=>	62902,
		20595	=>	62901,
		20596	=>	62899,
		20597	=>	62898,
		20598	=>	62897,
		20599	=>	62896,
		20600	=>	62894,
		20601	=>	62893,
		20602	=>	62892,
		20603	=>	62891,
		20604	=>	62890,
		20605	=>	62888,
		20606	=>	62887,
		20607	=>	62886,
		20608	=>	62885,
		20609	=>	62883,
		20610	=>	62882,
		20611	=>	62881,
		20612	=>	62880,
		20613	=>	62878,
		20614	=>	62877,
		20615	=>	62876,
		20616	=>	62875,
		20617	=>	62873,
		20618	=>	62872,
		20619	=>	62871,
		20620	=>	62870,
		20621	=>	62868,
		20622	=>	62867,
		20623	=>	62866,
		20624	=>	62865,
		20625	=>	62863,
		20626	=>	62862,
		20627	=>	62861,
		20628	=>	62860,
		20629	=>	62859,
		20630	=>	62857,
		20631	=>	62856,
		20632	=>	62855,
		20633	=>	62854,
		20634	=>	62852,
		20635	=>	62851,
		20636	=>	62850,
		20637	=>	62849,
		20638	=>	62847,
		20639	=>	62846,
		20640	=>	62845,
		20641	=>	62844,
		20642	=>	62842,
		20643	=>	62841,
		20644	=>	62840,
		20645	=>	62839,
		20646	=>	62837,
		20647	=>	62836,
		20648	=>	62835,
		20649	=>	62834,
		20650	=>	62832,
		20651	=>	62831,
		20652	=>	62830,
		20653	=>	62829,
		20654	=>	62827,
		20655	=>	62826,
		20656	=>	62825,
		20657	=>	62824,
		20658	=>	62822,
		20659	=>	62821,
		20660	=>	62820,
		20661	=>	62819,
		20662	=>	62817,
		20663	=>	62816,
		20664	=>	62815,
		20665	=>	62814,
		20666	=>	62812,
		20667	=>	62811,
		20668	=>	62810,
		20669	=>	62809,
		20670	=>	62807,
		20671	=>	62806,
		20672	=>	62805,
		20673	=>	62804,
		20674	=>	62802,
		20675	=>	62801,
		20676	=>	62800,
		20677	=>	62799,
		20678	=>	62797,
		20679	=>	62796,
		20680	=>	62795,
		20681	=>	62793,
		20682	=>	62792,
		20683	=>	62791,
		20684	=>	62790,
		20685	=>	62788,
		20686	=>	62787,
		20687	=>	62786,
		20688	=>	62785,
		20689	=>	62783,
		20690	=>	62782,
		20691	=>	62781,
		20692	=>	62780,
		20693	=>	62778,
		20694	=>	62777,
		20695	=>	62776,
		20696	=>	62775,
		20697	=>	62773,
		20698	=>	62772,
		20699	=>	62771,
		20700	=>	62770,
		20701	=>	62768,
		20702	=>	62767,
		20703	=>	62766,
		20704	=>	62764,
		20705	=>	62763,
		20706	=>	62762,
		20707	=>	62761,
		20708	=>	62759,
		20709	=>	62758,
		20710	=>	62757,
		20711	=>	62756,
		20712	=>	62754,
		20713	=>	62753,
		20714	=>	62752,
		20715	=>	62751,
		20716	=>	62749,
		20717	=>	62748,
		20718	=>	62747,
		20719	=>	62745,
		20720	=>	62744,
		20721	=>	62743,
		20722	=>	62742,
		20723	=>	62740,
		20724	=>	62739,
		20725	=>	62738,
		20726	=>	62737,
		20727	=>	62735,
		20728	=>	62734,
		20729	=>	62733,
		20730	=>	62732,
		20731	=>	62730,
		20732	=>	62729,
		20733	=>	62728,
		20734	=>	62726,
		20735	=>	62725,
		20736	=>	62724,
		20737	=>	62723,
		20738	=>	62721,
		20739	=>	62720,
		20740	=>	62719,
		20741	=>	62717,
		20742	=>	62716,
		20743	=>	62715,
		20744	=>	62714,
		20745	=>	62712,
		20746	=>	62711,
		20747	=>	62710,
		20748	=>	62709,
		20749	=>	62707,
		20750	=>	62706,
		20751	=>	62705,
		20752	=>	62703,
		20753	=>	62702,
		20754	=>	62701,
		20755	=>	62700,
		20756	=>	62698,
		20757	=>	62697,
		20758	=>	62696,
		20759	=>	62695,
		20760	=>	62693,
		20761	=>	62692,
		20762	=>	62691,
		20763	=>	62689,
		20764	=>	62688,
		20765	=>	62687,
		20766	=>	62686,
		20767	=>	62684,
		20768	=>	62683,
		20769	=>	62682,
		20770	=>	62680,
		20771	=>	62679,
		20772	=>	62678,
		20773	=>	62677,
		20774	=>	62675,
		20775	=>	62674,
		20776	=>	62673,
		20777	=>	62671,
		20778	=>	62670,
		20779	=>	62669,
		20780	=>	62668,
		20781	=>	62666,
		20782	=>	62665,
		20783	=>	62664,
		20784	=>	62662,
		20785	=>	62661,
		20786	=>	62660,
		20787	=>	62659,
		20788	=>	62657,
		20789	=>	62656,
		20790	=>	62655,
		20791	=>	62653,
		20792	=>	62652,
		20793	=>	62651,
		20794	=>	62650,
		20795	=>	62648,
		20796	=>	62647,
		20797	=>	62646,
		20798	=>	62644,
		20799	=>	62643,
		20800	=>	62642,
		20801	=>	62641,
		20802	=>	62639,
		20803	=>	62638,
		20804	=>	62637,
		20805	=>	62635,
		20806	=>	62634,
		20807	=>	62633,
		20808	=>	62631,
		20809	=>	62630,
		20810	=>	62629,
		20811	=>	62628,
		20812	=>	62626,
		20813	=>	62625,
		20814	=>	62624,
		20815	=>	62622,
		20816	=>	62621,
		20817	=>	62620,
		20818	=>	62619,
		20819	=>	62617,
		20820	=>	62616,
		20821	=>	62615,
		20822	=>	62613,
		20823	=>	62612,
		20824	=>	62611,
		20825	=>	62609,
		20826	=>	62608,
		20827	=>	62607,
		20828	=>	62606,
		20829	=>	62604,
		20830	=>	62603,
		20831	=>	62602,
		20832	=>	62600,
		20833	=>	62599,
		20834	=>	62598,
		20835	=>	62596,
		20836	=>	62595,
		20837	=>	62594,
		20838	=>	62593,
		20839	=>	62591,
		20840	=>	62590,
		20841	=>	62589,
		20842	=>	62587,
		20843	=>	62586,
		20844	=>	62585,
		20845	=>	62583,
		20846	=>	62582,
		20847	=>	62581,
		20848	=>	62580,
		20849	=>	62578,
		20850	=>	62577,
		20851	=>	62576,
		20852	=>	62574,
		20853	=>	62573,
		20854	=>	62572,
		20855	=>	62570,
		20856	=>	62569,
		20857	=>	62568,
		20858	=>	62567,
		20859	=>	62565,
		20860	=>	62564,
		20861	=>	62563,
		20862	=>	62561,
		20863	=>	62560,
		20864	=>	62559,
		20865	=>	62557,
		20866	=>	62556,
		20867	=>	62555,
		20868	=>	62553,
		20869	=>	62552,
		20870	=>	62551,
		20871	=>	62549,
		20872	=>	62548,
		20873	=>	62547,
		20874	=>	62546,
		20875	=>	62544,
		20876	=>	62543,
		20877	=>	62542,
		20878	=>	62540,
		20879	=>	62539,
		20880	=>	62538,
		20881	=>	62536,
		20882	=>	62535,
		20883	=>	62534,
		20884	=>	62532,
		20885	=>	62531,
		20886	=>	62530,
		20887	=>	62529,
		20888	=>	62527,
		20889	=>	62526,
		20890	=>	62525,
		20891	=>	62523,
		20892	=>	62522,
		20893	=>	62521,
		20894	=>	62519,
		20895	=>	62518,
		20896	=>	62517,
		20897	=>	62515,
		20898	=>	62514,
		20899	=>	62513,
		20900	=>	62511,
		20901	=>	62510,
		20902	=>	62509,
		20903	=>	62507,
		20904	=>	62506,
		20905	=>	62505,
		20906	=>	62503,
		20907	=>	62502,
		20908	=>	62501,
		20909	=>	62500,
		20910	=>	62498,
		20911	=>	62497,
		20912	=>	62496,
		20913	=>	62494,
		20914	=>	62493,
		20915	=>	62492,
		20916	=>	62490,
		20917	=>	62489,
		20918	=>	62488,
		20919	=>	62486,
		20920	=>	62485,
		20921	=>	62484,
		20922	=>	62482,
		20923	=>	62481,
		20924	=>	62480,
		20925	=>	62478,
		20926	=>	62477,
		20927	=>	62476,
		20928	=>	62474,
		20929	=>	62473,
		20930	=>	62472,
		20931	=>	62470,
		20932	=>	62469,
		20933	=>	62468,
		20934	=>	62466,
		20935	=>	62465,
		20936	=>	62464,
		20937	=>	62462,
		20938	=>	62461,
		20939	=>	62460,
		20940	=>	62458,
		20941	=>	62457,
		20942	=>	62456,
		20943	=>	62454,
		20944	=>	62453,
		20945	=>	62452,
		20946	=>	62450,
		20947	=>	62449,
		20948	=>	62448,
		20949	=>	62446,
		20950	=>	62445,
		20951	=>	62444,
		20952	=>	62442,
		20953	=>	62441,
		20954	=>	62440,
		20955	=>	62438,
		20956	=>	62437,
		20957	=>	62436,
		20958	=>	62434,
		20959	=>	62433,
		20960	=>	62432,
		20961	=>	62430,
		20962	=>	62429,
		20963	=>	62428,
		20964	=>	62426,
		20965	=>	62425,
		20966	=>	62424,
		20967	=>	62422,
		20968	=>	62421,
		20969	=>	62420,
		20970	=>	62418,
		20971	=>	62417,
		20972	=>	62416,
		20973	=>	62414,
		20974	=>	62413,
		20975	=>	62412,
		20976	=>	62410,
		20977	=>	62409,
		20978	=>	62408,
		20979	=>	62406,
		20980	=>	62405,
		20981	=>	62404,
		20982	=>	62402,
		20983	=>	62401,
		20984	=>	62400,
		20985	=>	62398,
		20986	=>	62397,
		20987	=>	62396,
		20988	=>	62394,
		20989	=>	62393,
		20990	=>	62392,
		20991	=>	62390,
		20992	=>	62389,
		20993	=>	62388,
		20994	=>	62386,
		20995	=>	62385,
		20996	=>	62384,
		20997	=>	62382,
		20998	=>	62381,
		20999	=>	62380,
		21000	=>	62378,
		21001	=>	62377,
		21002	=>	62376,
		21003	=>	62374,
		21004	=>	62373,
		21005	=>	62371,
		21006	=>	62370,
		21007	=>	62369,
		21008	=>	62367,
		21009	=>	62366,
		21010	=>	62365,
		21011	=>	62363,
		21012	=>	62362,
		21013	=>	62361,
		21014	=>	62359,
		21015	=>	62358,
		21016	=>	62357,
		21017	=>	62355,
		21018	=>	62354,
		21019	=>	62353,
		21020	=>	62351,
		21021	=>	62350,
		21022	=>	62349,
		21023	=>	62347,
		21024	=>	62346,
		21025	=>	62344,
		21026	=>	62343,
		21027	=>	62342,
		21028	=>	62340,
		21029	=>	62339,
		21030	=>	62338,
		21031	=>	62336,
		21032	=>	62335,
		21033	=>	62334,
		21034	=>	62332,
		21035	=>	62331,
		21036	=>	62330,
		21037	=>	62328,
		21038	=>	62327,
		21039	=>	62326,
		21040	=>	62324,
		21041	=>	62323,
		21042	=>	62321,
		21043	=>	62320,
		21044	=>	62319,
		21045	=>	62317,
		21046	=>	62316,
		21047	=>	62315,
		21048	=>	62313,
		21049	=>	62312,
		21050	=>	62311,
		21051	=>	62309,
		21052	=>	62308,
		21053	=>	62307,
		21054	=>	62305,
		21055	=>	62304,
		21056	=>	62302,
		21057	=>	62301,
		21058	=>	62300,
		21059	=>	62298,
		21060	=>	62297,
		21061	=>	62296,
		21062	=>	62294,
		21063	=>	62293,
		21064	=>	62292,
		21065	=>	62290,
		21066	=>	62289,
		21067	=>	62287,
		21068	=>	62286,
		21069	=>	62285,
		21070	=>	62283,
		21071	=>	62282,
		21072	=>	62281,
		21073	=>	62279,
		21074	=>	62278,
		21075	=>	62277,
		21076	=>	62275,
		21077	=>	62274,
		21078	=>	62272,
		21079	=>	62271,
		21080	=>	62270,
		21081	=>	62268,
		21082	=>	62267,
		21083	=>	62266,
		21084	=>	62264,
		21085	=>	62263,
		21086	=>	62262,
		21087	=>	62260,
		21088	=>	62259,
		21089	=>	62257,
		21090	=>	62256,
		21091	=>	62255,
		21092	=>	62253,
		21093	=>	62252,
		21094	=>	62251,
		21095	=>	62249,
		21096	=>	62248,
		21097	=>	62246,
		21098	=>	62245,
		21099	=>	62244,
		21100	=>	62242,
		21101	=>	62241,
		21102	=>	62240,
		21103	=>	62238,
		21104	=>	62237,
		21105	=>	62235,
		21106	=>	62234,
		21107	=>	62233,
		21108	=>	62231,
		21109	=>	62230,
		21110	=>	62229,
		21111	=>	62227,
		21112	=>	62226,
		21113	=>	62224,
		21114	=>	62223,
		21115	=>	62222,
		21116	=>	62220,
		21117	=>	62219,
		21118	=>	62218,
		21119	=>	62216,
		21120	=>	62215,
		21121	=>	62213,
		21122	=>	62212,
		21123	=>	62211,
		21124	=>	62209,
		21125	=>	62208,
		21126	=>	62207,
		21127	=>	62205,
		21128	=>	62204,
		21129	=>	62202,
		21130	=>	62201,
		21131	=>	62200,
		21132	=>	62198,
		21133	=>	62197,
		21134	=>	62195,
		21135	=>	62194,
		21136	=>	62193,
		21137	=>	62191,
		21138	=>	62190,
		21139	=>	62189,
		21140	=>	62187,
		21141	=>	62186,
		21142	=>	62184,
		21143	=>	62183,
		21144	=>	62182,
		21145	=>	62180,
		21146	=>	62179,
		21147	=>	62178,
		21148	=>	62176,
		21149	=>	62175,
		21150	=>	62173,
		21151	=>	62172,
		21152	=>	62171,
		21153	=>	62169,
		21154	=>	62168,
		21155	=>	62166,
		21156	=>	62165,
		21157	=>	62164,
		21158	=>	62162,
		21159	=>	62161,
		21160	=>	62159,
		21161	=>	62158,
		21162	=>	62157,
		21163	=>	62155,
		21164	=>	62154,
		21165	=>	62153,
		21166	=>	62151,
		21167	=>	62150,
		21168	=>	62148,
		21169	=>	62147,
		21170	=>	62146,
		21171	=>	62144,
		21172	=>	62143,
		21173	=>	62141,
		21174	=>	62140,
		21175	=>	62139,
		21176	=>	62137,
		21177	=>	62136,
		21178	=>	62134,
		21179	=>	62133,
		21180	=>	62132,
		21181	=>	62130,
		21182	=>	62129,
		21183	=>	62127,
		21184	=>	62126,
		21185	=>	62125,
		21186	=>	62123,
		21187	=>	62122,
		21188	=>	62120,
		21189	=>	62119,
		21190	=>	62118,
		21191	=>	62116,
		21192	=>	62115,
		21193	=>	62114,
		21194	=>	62112,
		21195	=>	62111,
		21196	=>	62109,
		21197	=>	62108,
		21198	=>	62107,
		21199	=>	62105,
		21200	=>	62104,
		21201	=>	62102,
		21202	=>	62101,
		21203	=>	62100,
		21204	=>	62098,
		21205	=>	62097,
		21206	=>	62095,
		21207	=>	62094,
		21208	=>	62093,
		21209	=>	62091,
		21210	=>	62090,
		21211	=>	62088,
		21212	=>	62087,
		21213	=>	62085,
		21214	=>	62084,
		21215	=>	62083,
		21216	=>	62081,
		21217	=>	62080,
		21218	=>	62078,
		21219	=>	62077,
		21220	=>	62076,
		21221	=>	62074,
		21222	=>	62073,
		21223	=>	62071,
		21224	=>	62070,
		21225	=>	62069,
		21226	=>	62067,
		21227	=>	62066,
		21228	=>	62064,
		21229	=>	62063,
		21230	=>	62062,
		21231	=>	62060,
		21232	=>	62059,
		21233	=>	62057,
		21234	=>	62056,
		21235	=>	62055,
		21236	=>	62053,
		21237	=>	62052,
		21238	=>	62050,
		21239	=>	62049,
		21240	=>	62048,
		21241	=>	62046,
		21242	=>	62045,
		21243	=>	62043,
		21244	=>	62042,
		21245	=>	62040,
		21246	=>	62039,
		21247	=>	62038,
		21248	=>	62036,
		21249	=>	62035,
		21250	=>	62033,
		21251	=>	62032,
		21252	=>	62031,
		21253	=>	62029,
		21254	=>	62028,
		21255	=>	62026,
		21256	=>	62025,
		21257	=>	62024,
		21258	=>	62022,
		21259	=>	62021,
		21260	=>	62019,
		21261	=>	62018,
		21262	=>	62016,
		21263	=>	62015,
		21264	=>	62014,
		21265	=>	62012,
		21266	=>	62011,
		21267	=>	62009,
		21268	=>	62008,
		21269	=>	62007,
		21270	=>	62005,
		21271	=>	62004,
		21272	=>	62002,
		21273	=>	62001,
		21274	=>	61999,
		21275	=>	61998,
		21276	=>	61997,
		21277	=>	61995,
		21278	=>	61994,
		21279	=>	61992,
		21280	=>	61991,
		21281	=>	61989,
		21282	=>	61988,
		21283	=>	61987,
		21284	=>	61985,
		21285	=>	61984,
		21286	=>	61982,
		21287	=>	61981,
		21288	=>	61980,
		21289	=>	61978,
		21290	=>	61977,
		21291	=>	61975,
		21292	=>	61974,
		21293	=>	61972,
		21294	=>	61971,
		21295	=>	61970,
		21296	=>	61968,
		21297	=>	61967,
		21298	=>	61965,
		21299	=>	61964,
		21300	=>	61962,
		21301	=>	61961,
		21302	=>	61960,
		21303	=>	61958,
		21304	=>	61957,
		21305	=>	61955,
		21306	=>	61954,
		21307	=>	61952,
		21308	=>	61951,
		21309	=>	61950,
		21310	=>	61948,
		21311	=>	61947,
		21312	=>	61945,
		21313	=>	61944,
		21314	=>	61942,
		21315	=>	61941,
		21316	=>	61940,
		21317	=>	61938,
		21318	=>	61937,
		21319	=>	61935,
		21320	=>	61934,
		21321	=>	61932,
		21322	=>	61931,
		21323	=>	61930,
		21324	=>	61928,
		21325	=>	61927,
		21326	=>	61925,
		21327	=>	61924,
		21328	=>	61922,
		21329	=>	61921,
		21330	=>	61920,
		21331	=>	61918,
		21332	=>	61917,
		21333	=>	61915,
		21334	=>	61914,
		21335	=>	61912,
		21336	=>	61911,
		21337	=>	61909,
		21338	=>	61908,
		21339	=>	61907,
		21340	=>	61905,
		21341	=>	61904,
		21342	=>	61902,
		21343	=>	61901,
		21344	=>	61899,
		21345	=>	61898,
		21346	=>	61897,
		21347	=>	61895,
		21348	=>	61894,
		21349	=>	61892,
		21350	=>	61891,
		21351	=>	61889,
		21352	=>	61888,
		21353	=>	61886,
		21354	=>	61885,
		21355	=>	61884,
		21356	=>	61882,
		21357	=>	61881,
		21358	=>	61879,
		21359	=>	61878,
		21360	=>	61876,
		21361	=>	61875,
		21362	=>	61873,
		21363	=>	61872,
		21364	=>	61871,
		21365	=>	61869,
		21366	=>	61868,
		21367	=>	61866,
		21368	=>	61865,
		21369	=>	61863,
		21370	=>	61862,
		21371	=>	61860,
		21372	=>	61859,
		21373	=>	61858,
		21374	=>	61856,
		21375	=>	61855,
		21376	=>	61853,
		21377	=>	61852,
		21378	=>	61850,
		21379	=>	61849,
		21380	=>	61847,
		21381	=>	61846,
		21382	=>	61845,
		21383	=>	61843,
		21384	=>	61842,
		21385	=>	61840,
		21386	=>	61839,
		21387	=>	61837,
		21388	=>	61836,
		21389	=>	61834,
		21390	=>	61833,
		21391	=>	61831,
		21392	=>	61830,
		21393	=>	61829,
		21394	=>	61827,
		21395	=>	61826,
		21396	=>	61824,
		21397	=>	61823,
		21398	=>	61821,
		21399	=>	61820,
		21400	=>	61818,
		21401	=>	61817,
		21402	=>	61816,
		21403	=>	61814,
		21404	=>	61813,
		21405	=>	61811,
		21406	=>	61810,
		21407	=>	61808,
		21408	=>	61807,
		21409	=>	61805,
		21410	=>	61804,
		21411	=>	61802,
		21412	=>	61801,
		21413	=>	61800,
		21414	=>	61798,
		21415	=>	61797,
		21416	=>	61795,
		21417	=>	61794,
		21418	=>	61792,
		21419	=>	61791,
		21420	=>	61789,
		21421	=>	61788,
		21422	=>	61786,
		21423	=>	61785,
		21424	=>	61783,
		21425	=>	61782,
		21426	=>	61781,
		21427	=>	61779,
		21428	=>	61778,
		21429	=>	61776,
		21430	=>	61775,
		21431	=>	61773,
		21432	=>	61772,
		21433	=>	61770,
		21434	=>	61769,
		21435	=>	61767,
		21436	=>	61766,
		21437	=>	61764,
		21438	=>	61763,
		21439	=>	61762,
		21440	=>	61760,
		21441	=>	61759,
		21442	=>	61757,
		21443	=>	61756,
		21444	=>	61754,
		21445	=>	61753,
		21446	=>	61751,
		21447	=>	61750,
		21448	=>	61748,
		21449	=>	61747,
		21450	=>	61745,
		21451	=>	61744,
		21452	=>	61743,
		21453	=>	61741,
		21454	=>	61740,
		21455	=>	61738,
		21456	=>	61737,
		21457	=>	61735,
		21458	=>	61734,
		21459	=>	61732,
		21460	=>	61731,
		21461	=>	61729,
		21462	=>	61728,
		21463	=>	61726,
		21464	=>	61725,
		21465	=>	61723,
		21466	=>	61722,
		21467	=>	61720,
		21468	=>	61719,
		21469	=>	61718,
		21470	=>	61716,
		21471	=>	61715,
		21472	=>	61713,
		21473	=>	61712,
		21474	=>	61710,
		21475	=>	61709,
		21476	=>	61707,
		21477	=>	61706,
		21478	=>	61704,
		21479	=>	61703,
		21480	=>	61701,
		21481	=>	61700,
		21482	=>	61698,
		21483	=>	61697,
		21484	=>	61695,
		21485	=>	61694,
		21486	=>	61692,
		21487	=>	61691,
		21488	=>	61690,
		21489	=>	61688,
		21490	=>	61687,
		21491	=>	61685,
		21492	=>	61684,
		21493	=>	61682,
		21494	=>	61681,
		21495	=>	61679,
		21496	=>	61678,
		21497	=>	61676,
		21498	=>	61675,
		21499	=>	61673,
		21500	=>	61672,
		21501	=>	61670,
		21502	=>	61669,
		21503	=>	61667,
		21504	=>	61666,
		21505	=>	61664,
		21506	=>	61663,
		21507	=>	61661,
		21508	=>	61660,
		21509	=>	61658,
		21510	=>	61657,
		21511	=>	61655,
		21512	=>	61654,
		21513	=>	61653,
		21514	=>	61651,
		21515	=>	61650,
		21516	=>	61648,
		21517	=>	61647,
		21518	=>	61645,
		21519	=>	61644,
		21520	=>	61642,
		21521	=>	61641,
		21522	=>	61639,
		21523	=>	61638,
		21524	=>	61636,
		21525	=>	61635,
		21526	=>	61633,
		21527	=>	61632,
		21528	=>	61630,
		21529	=>	61629,
		21530	=>	61627,
		21531	=>	61626,
		21532	=>	61624,
		21533	=>	61623,
		21534	=>	61621,
		21535	=>	61620,
		21536	=>	61618,
		21537	=>	61617,
		21538	=>	61615,
		21539	=>	61614,
		21540	=>	61612,
		21541	=>	61611,
		21542	=>	61609,
		21543	=>	61608,
		21544	=>	61606,
		21545	=>	61605,
		21546	=>	61603,
		21547	=>	61602,
		21548	=>	61600,
		21549	=>	61599,
		21550	=>	61597,
		21551	=>	61596,
		21552	=>	61594,
		21553	=>	61593,
		21554	=>	61591,
		21555	=>	61590,
		21556	=>	61588,
		21557	=>	61587,
		21558	=>	61585,
		21559	=>	61584,
		21560	=>	61583,
		21561	=>	61581,
		21562	=>	61580,
		21563	=>	61578,
		21564	=>	61577,
		21565	=>	61575,
		21566	=>	61574,
		21567	=>	61572,
		21568	=>	61571,
		21569	=>	61569,
		21570	=>	61568,
		21571	=>	61566,
		21572	=>	61565,
		21573	=>	61563,
		21574	=>	61562,
		21575	=>	61560,
		21576	=>	61559,
		21577	=>	61557,
		21578	=>	61556,
		21579	=>	61554,
		21580	=>	61553,
		21581	=>	61551,
		21582	=>	61550,
		21583	=>	61548,
		21584	=>	61547,
		21585	=>	61545,
		21586	=>	61544,
		21587	=>	61542,
		21588	=>	61541,
		21589	=>	61539,
		21590	=>	61538,
		21591	=>	61536,
		21592	=>	61535,
		21593	=>	61533,
		21594	=>	61531,
		21595	=>	61530,
		21596	=>	61528,
		21597	=>	61527,
		21598	=>	61525,
		21599	=>	61524,
		21600	=>	61522,
		21601	=>	61521,
		21602	=>	61519,
		21603	=>	61518,
		21604	=>	61516,
		21605	=>	61515,
		21606	=>	61513,
		21607	=>	61512,
		21608	=>	61510,
		21609	=>	61509,
		21610	=>	61507,
		21611	=>	61506,
		21612	=>	61504,
		21613	=>	61503,
		21614	=>	61501,
		21615	=>	61500,
		21616	=>	61498,
		21617	=>	61497,
		21618	=>	61495,
		21619	=>	61494,
		21620	=>	61492,
		21621	=>	61491,
		21622	=>	61489,
		21623	=>	61488,
		21624	=>	61486,
		21625	=>	61485,
		21626	=>	61483,
		21627	=>	61482,
		21628	=>	61480,
		21629	=>	61479,
		21630	=>	61477,
		21631	=>	61476,
		21632	=>	61474,
		21633	=>	61473,
		21634	=>	61471,
		21635	=>	61470,
		21636	=>	61468,
		21637	=>	61467,
		21638	=>	61465,
		21639	=>	61464,
		21640	=>	61462,
		21641	=>	61460,
		21642	=>	61459,
		21643	=>	61457,
		21644	=>	61456,
		21645	=>	61454,
		21646	=>	61453,
		21647	=>	61451,
		21648	=>	61450,
		21649	=>	61448,
		21650	=>	61447,
		21651	=>	61445,
		21652	=>	61444,
		21653	=>	61442,
		21654	=>	61441,
		21655	=>	61439,
		21656	=>	61438,
		21657	=>	61436,
		21658	=>	61435,
		21659	=>	61433,
		21660	=>	61432,
		21661	=>	61430,
		21662	=>	61429,
		21663	=>	61427,
		21664	=>	61426,
		21665	=>	61424,
		21666	=>	61422,
		21667	=>	61421,
		21668	=>	61419,
		21669	=>	61418,
		21670	=>	61416,
		21671	=>	61415,
		21672	=>	61413,
		21673	=>	61412,
		21674	=>	61410,
		21675	=>	61409,
		21676	=>	61407,
		21677	=>	61406,
		21678	=>	61404,
		21679	=>	61403,
		21680	=>	61401,
		21681	=>	61400,
		21682	=>	61398,
		21683	=>	61397,
		21684	=>	61395,
		21685	=>	61393,
		21686	=>	61392,
		21687	=>	61390,
		21688	=>	61389,
		21689	=>	61387,
		21690	=>	61386,
		21691	=>	61384,
		21692	=>	61383,
		21693	=>	61381,
		21694	=>	61380,
		21695	=>	61378,
		21696	=>	61377,
		21697	=>	61375,
		21698	=>	61374,
		21699	=>	61372,
		21700	=>	61371,
		21701	=>	61369,
		21702	=>	61367,
		21703	=>	61366,
		21704	=>	61364,
		21705	=>	61363,
		21706	=>	61361,
		21707	=>	61360,
		21708	=>	61358,
		21709	=>	61357,
		21710	=>	61355,
		21711	=>	61354,
		21712	=>	61352,
		21713	=>	61351,
		21714	=>	61349,
		21715	=>	61347,
		21716	=>	61346,
		21717	=>	61344,
		21718	=>	61343,
		21719	=>	61341,
		21720	=>	61340,
		21721	=>	61338,
		21722	=>	61337,
		21723	=>	61335,
		21724	=>	61334,
		21725	=>	61332,
		21726	=>	61331,
		21727	=>	61329,
		21728	=>	61327,
		21729	=>	61326,
		21730	=>	61324,
		21731	=>	61323,
		21732	=>	61321,
		21733	=>	61320,
		21734	=>	61318,
		21735	=>	61317,
		21736	=>	61315,
		21737	=>	61314,
		21738	=>	61312,
		21739	=>	61311,
		21740	=>	61309,
		21741	=>	61307,
		21742	=>	61306,
		21743	=>	61304,
		21744	=>	61303,
		21745	=>	61301,
		21746	=>	61300,
		21747	=>	61298,
		21748	=>	61297,
		21749	=>	61295,
		21750	=>	61294,
		21751	=>	61292,
		21752	=>	61290,
		21753	=>	61289,
		21754	=>	61287,
		21755	=>	61286,
		21756	=>	61284,
		21757	=>	61283,
		21758	=>	61281,
		21759	=>	61280,
		21760	=>	61278,
		21761	=>	61277,
		21762	=>	61275,
		21763	=>	61273,
		21764	=>	61272,
		21765	=>	61270,
		21766	=>	61269,
		21767	=>	61267,
		21768	=>	61266,
		21769	=>	61264,
		21770	=>	61263,
		21771	=>	61261,
		21772	=>	61259,
		21773	=>	61258,
		21774	=>	61256,
		21775	=>	61255,
		21776	=>	61253,
		21777	=>	61252,
		21778	=>	61250,
		21779	=>	61249,
		21780	=>	61247,
		21781	=>	61246,
		21782	=>	61244,
		21783	=>	61242,
		21784	=>	61241,
		21785	=>	61239,
		21786	=>	61238,
		21787	=>	61236,
		21788	=>	61235,
		21789	=>	61233,
		21790	=>	61232,
		21791	=>	61230,
		21792	=>	61228,
		21793	=>	61227,
		21794	=>	61225,
		21795	=>	61224,
		21796	=>	61222,
		21797	=>	61221,
		21798	=>	61219,
		21799	=>	61217,
		21800	=>	61216,
		21801	=>	61214,
		21802	=>	61213,
		21803	=>	61211,
		21804	=>	61210,
		21805	=>	61208,
		21806	=>	61207,
		21807	=>	61205,
		21808	=>	61203,
		21809	=>	61202,
		21810	=>	61200,
		21811	=>	61199,
		21812	=>	61197,
		21813	=>	61196,
		21814	=>	61194,
		21815	=>	61193,
		21816	=>	61191,
		21817	=>	61189,
		21818	=>	61188,
		21819	=>	61186,
		21820	=>	61185,
		21821	=>	61183,
		21822	=>	61182,
		21823	=>	61180,
		21824	=>	61178,
		21825	=>	61177,
		21826	=>	61175,
		21827	=>	61174,
		21828	=>	61172,
		21829	=>	61171,
		21830	=>	61169,
		21831	=>	61167,
		21832	=>	61166,
		21833	=>	61164,
		21834	=>	61163,
		21835	=>	61161,
		21836	=>	61160,
		21837	=>	61158,
		21838	=>	61156,
		21839	=>	61155,
		21840	=>	61153,
		21841	=>	61152,
		21842	=>	61150,
		21843	=>	61149,
		21844	=>	61147,
		21845	=>	61146,
		21846	=>	61144,
		21847	=>	61142,
		21848	=>	61141,
		21849	=>	61139,
		21850	=>	61138,
		21851	=>	61136,
		21852	=>	61135,
		21853	=>	61133,
		21854	=>	61131,
		21855	=>	61130,
		21856	=>	61128,
		21857	=>	61127,
		21858	=>	61125,
		21859	=>	61123,
		21860	=>	61122,
		21861	=>	61120,
		21862	=>	61119,
		21863	=>	61117,
		21864	=>	61116,
		21865	=>	61114,
		21866	=>	61112,
		21867	=>	61111,
		21868	=>	61109,
		21869	=>	61108,
		21870	=>	61106,
		21871	=>	61105,
		21872	=>	61103,
		21873	=>	61101,
		21874	=>	61100,
		21875	=>	61098,
		21876	=>	61097,
		21877	=>	61095,
		21878	=>	61094,
		21879	=>	61092,
		21880	=>	61090,
		21881	=>	61089,
		21882	=>	61087,
		21883	=>	61086,
		21884	=>	61084,
		21885	=>	61082,
		21886	=>	61081,
		21887	=>	61079,
		21888	=>	61078,
		21889	=>	61076,
		21890	=>	61075,
		21891	=>	61073,
		21892	=>	61071,
		21893	=>	61070,
		21894	=>	61068,
		21895	=>	61067,
		21896	=>	61065,
		21897	=>	61063,
		21898	=>	61062,
		21899	=>	61060,
		21900	=>	61059,
		21901	=>	61057,
		21902	=>	61056,
		21903	=>	61054,
		21904	=>	61052,
		21905	=>	61051,
		21906	=>	61049,
		21907	=>	61048,
		21908	=>	61046,
		21909	=>	61044,
		21910	=>	61043,
		21911	=>	61041,
		21912	=>	61040,
		21913	=>	61038,
		21914	=>	61037,
		21915	=>	61035,
		21916	=>	61033,
		21917	=>	61032,
		21918	=>	61030,
		21919	=>	61029,
		21920	=>	61027,
		21921	=>	61025,
		21922	=>	61024,
		21923	=>	61022,
		21924	=>	61021,
		21925	=>	61019,
		21926	=>	61017,
		21927	=>	61016,
		21928	=>	61014,
		21929	=>	61013,
		21930	=>	61011,
		21931	=>	61009,
		21932	=>	61008,
		21933	=>	61006,
		21934	=>	61005,
		21935	=>	61003,
		21936	=>	61002,
		21937	=>	61000,
		21938	=>	60998,
		21939	=>	60997,
		21940	=>	60995,
		21941	=>	60994,
		21942	=>	60992,
		21943	=>	60990,
		21944	=>	60989,
		21945	=>	60987,
		21946	=>	60986,
		21947	=>	60984,
		21948	=>	60982,
		21949	=>	60981,
		21950	=>	60979,
		21951	=>	60978,
		21952	=>	60976,
		21953	=>	60974,
		21954	=>	60973,
		21955	=>	60971,
		21956	=>	60970,
		21957	=>	60968,
		21958	=>	60966,
		21959	=>	60965,
		21960	=>	60963,
		21961	=>	60962,
		21962	=>	60960,
		21963	=>	60958,
		21964	=>	60957,
		21965	=>	60955,
		21966	=>	60954,
		21967	=>	60952,
		21968	=>	60950,
		21969	=>	60949,
		21970	=>	60947,
		21971	=>	60946,
		21972	=>	60944,
		21973	=>	60942,
		21974	=>	60941,
		21975	=>	60939,
		21976	=>	60938,
		21977	=>	60936,
		21978	=>	60934,
		21979	=>	60933,
		21980	=>	60931,
		21981	=>	60929,
		21982	=>	60928,
		21983	=>	60926,
		21984	=>	60925,
		21985	=>	60923,
		21986	=>	60921,
		21987	=>	60920,
		21988	=>	60918,
		21989	=>	60917,
		21990	=>	60915,
		21991	=>	60913,
		21992	=>	60912,
		21993	=>	60910,
		21994	=>	60909,
		21995	=>	60907,
		21996	=>	60905,
		21997	=>	60904,
		21998	=>	60902,
		21999	=>	60901,
		22000	=>	60899,
		22001	=>	60897,
		22002	=>	60896,
		22003	=>	60894,
		22004	=>	60892,
		22005	=>	60891,
		22006	=>	60889,
		22007	=>	60888,
		22008	=>	60886,
		22009	=>	60884,
		22010	=>	60883,
		22011	=>	60881,
		22012	=>	60880,
		22013	=>	60878,
		22014	=>	60876,
		22015	=>	60875,
		22016	=>	60873,
		22017	=>	60872,
		22018	=>	60870,
		22019	=>	60868,
		22020	=>	60867,
		22021	=>	60865,
		22022	=>	60863,
		22023	=>	60862,
		22024	=>	60860,
		22025	=>	60859,
		22026	=>	60857,
		22027	=>	60855,
		22028	=>	60854,
		22029	=>	60852,
		22030	=>	60850,
		22031	=>	60849,
		22032	=>	60847,
		22033	=>	60846,
		22034	=>	60844,
		22035	=>	60842,
		22036	=>	60841,
		22037	=>	60839,
		22038	=>	60838,
		22039	=>	60836,
		22040	=>	60834,
		22041	=>	60833,
		22042	=>	60831,
		22043	=>	60829,
		22044	=>	60828,
		22045	=>	60826,
		22046	=>	60825,
		22047	=>	60823,
		22048	=>	60821,
		22049	=>	60820,
		22050	=>	60818,
		22051	=>	60816,
		22052	=>	60815,
		22053	=>	60813,
		22054	=>	60812,
		22055	=>	60810,
		22056	=>	60808,
		22057	=>	60807,
		22058	=>	60805,
		22059	=>	60803,
		22060	=>	60802,
		22061	=>	60800,
		22062	=>	60799,
		22063	=>	60797,
		22064	=>	60795,
		22065	=>	60794,
		22066	=>	60792,
		22067	=>	60790,
		22068	=>	60789,
		22069	=>	60787,
		22070	=>	60786,
		22071	=>	60784,
		22072	=>	60782,
		22073	=>	60781,
		22074	=>	60779,
		22075	=>	60777,
		22076	=>	60776,
		22077	=>	60774,
		22078	=>	60772,
		22079	=>	60771,
		22080	=>	60769,
		22081	=>	60768,
		22082	=>	60766,
		22083	=>	60764,
		22084	=>	60763,
		22085	=>	60761,
		22086	=>	60759,
		22087	=>	60758,
		22088	=>	60756,
		22089	=>	60755,
		22090	=>	60753,
		22091	=>	60751,
		22092	=>	60750,
		22093	=>	60748,
		22094	=>	60746,
		22095	=>	60745,
		22096	=>	60743,
		22097	=>	60741,
		22098	=>	60740,
		22099	=>	60738,
		22100	=>	60737,
		22101	=>	60735,
		22102	=>	60733,
		22103	=>	60732,
		22104	=>	60730,
		22105	=>	60728,
		22106	=>	60727,
		22107	=>	60725,
		22108	=>	60723,
		22109	=>	60722,
		22110	=>	60720,
		22111	=>	60719,
		22112	=>	60717,
		22113	=>	60715,
		22114	=>	60714,
		22115	=>	60712,
		22116	=>	60710,
		22117	=>	60709,
		22118	=>	60707,
		22119	=>	60705,
		22120	=>	60704,
		22121	=>	60702,
		22122	=>	60700,
		22123	=>	60699,
		22124	=>	60697,
		22125	=>	60696,
		22126	=>	60694,
		22127	=>	60692,
		22128	=>	60691,
		22129	=>	60689,
		22130	=>	60687,
		22131	=>	60686,
		22132	=>	60684,
		22133	=>	60682,
		22134	=>	60681,
		22135	=>	60679,
		22136	=>	60677,
		22137	=>	60676,
		22138	=>	60674,
		22139	=>	60673,
		22140	=>	60671,
		22141	=>	60669,
		22142	=>	60668,
		22143	=>	60666,
		22144	=>	60664,
		22145	=>	60663,
		22146	=>	60661,
		22147	=>	60659,
		22148	=>	60658,
		22149	=>	60656,
		22150	=>	60654,
		22151	=>	60653,
		22152	=>	60651,
		22153	=>	60649,
		22154	=>	60648,
		22155	=>	60646,
		22156	=>	60644,
		22157	=>	60643,
		22158	=>	60641,
		22159	=>	60640,
		22160	=>	60638,
		22161	=>	60636,
		22162	=>	60635,
		22163	=>	60633,
		22164	=>	60631,
		22165	=>	60630,
		22166	=>	60628,
		22167	=>	60626,
		22168	=>	60625,
		22169	=>	60623,
		22170	=>	60621,
		22171	=>	60620,
		22172	=>	60618,
		22173	=>	60616,
		22174	=>	60615,
		22175	=>	60613,
		22176	=>	60611,
		22177	=>	60610,
		22178	=>	60608,
		22179	=>	60606,
		22180	=>	60605,
		22181	=>	60603,
		22182	=>	60601,
		22183	=>	60600,
		22184	=>	60598,
		22185	=>	60596,
		22186	=>	60595,
		22187	=>	60593,
		22188	=>	60592,
		22189	=>	60590,
		22190	=>	60588,
		22191	=>	60587,
		22192	=>	60585,
		22193	=>	60583,
		22194	=>	60582,
		22195	=>	60580,
		22196	=>	60578,
		22197	=>	60577,
		22198	=>	60575,
		22199	=>	60573,
		22200	=>	60572,
		22201	=>	60570,
		22202	=>	60568,
		22203	=>	60567,
		22204	=>	60565,
		22205	=>	60563,
		22206	=>	60562,
		22207	=>	60560,
		22208	=>	60558,
		22209	=>	60557,
		22210	=>	60555,
		22211	=>	60553,
		22212	=>	60552,
		22213	=>	60550,
		22214	=>	60548,
		22215	=>	60547,
		22216	=>	60545,
		22217	=>	60543,
		22218	=>	60542,
		22219	=>	60540,
		22220	=>	60538,
		22221	=>	60537,
		22222	=>	60535,
		22223	=>	60533,
		22224	=>	60532,
		22225	=>	60530,
		22226	=>	60528,
		22227	=>	60527,
		22228	=>	60525,
		22229	=>	60523,
		22230	=>	60522,
		22231	=>	60520,
		22232	=>	60518,
		22233	=>	60517,
		22234	=>	60515,
		22235	=>	60513,
		22236	=>	60512,
		22237	=>	60510,
		22238	=>	60508,
		22239	=>	60507,
		22240	=>	60505,
		22241	=>	60503,
		22242	=>	60502,
		22243	=>	60500,
		22244	=>	60498,
		22245	=>	60497,
		22246	=>	60495,
		22247	=>	60493,
		22248	=>	60492,
		22249	=>	60490,
		22250	=>	60488,
		22251	=>	60486,
		22252	=>	60485,
		22253	=>	60483,
		22254	=>	60481,
		22255	=>	60480,
		22256	=>	60478,
		22257	=>	60476,
		22258	=>	60475,
		22259	=>	60473,
		22260	=>	60471,
		22261	=>	60470,
		22262	=>	60468,
		22263	=>	60466,
		22264	=>	60465,
		22265	=>	60463,
		22266	=>	60461,
		22267	=>	60460,
		22268	=>	60458,
		22269	=>	60456,
		22270	=>	60455,
		22271	=>	60453,
		22272	=>	60451,
		22273	=>	60450,
		22274	=>	60448,
		22275	=>	60446,
		22276	=>	60445,
		22277	=>	60443,
		22278	=>	60441,
		22279	=>	60439,
		22280	=>	60438,
		22281	=>	60436,
		22282	=>	60434,
		22283	=>	60433,
		22284	=>	60431,
		22285	=>	60429,
		22286	=>	60428,
		22287	=>	60426,
		22288	=>	60424,
		22289	=>	60423,
		22290	=>	60421,
		22291	=>	60419,
		22292	=>	60418,
		22293	=>	60416,
		22294	=>	60414,
		22295	=>	60413,
		22296	=>	60411,
		22297	=>	60409,
		22298	=>	60407,
		22299	=>	60406,
		22300	=>	60404,
		22301	=>	60402,
		22302	=>	60401,
		22303	=>	60399,
		22304	=>	60397,
		22305	=>	60396,
		22306	=>	60394,
		22307	=>	60392,
		22308	=>	60391,
		22309	=>	60389,
		22310	=>	60387,
		22311	=>	60385,
		22312	=>	60384,
		22313	=>	60382,
		22314	=>	60380,
		22315	=>	60379,
		22316	=>	60377,
		22317	=>	60375,
		22318	=>	60374,
		22319	=>	60372,
		22320	=>	60370,
		22321	=>	60369,
		22322	=>	60367,
		22323	=>	60365,
		22324	=>	60363,
		22325	=>	60362,
		22326	=>	60360,
		22327	=>	60358,
		22328	=>	60357,
		22329	=>	60355,
		22330	=>	60353,
		22331	=>	60352,
		22332	=>	60350,
		22333	=>	60348,
		22334	=>	60347,
		22335	=>	60345,
		22336	=>	60343,
		22337	=>	60341,
		22338	=>	60340,
		22339	=>	60338,
		22340	=>	60336,
		22341	=>	60335,
		22342	=>	60333,
		22343	=>	60331,
		22344	=>	60330,
		22345	=>	60328,
		22346	=>	60326,
		22347	=>	60324,
		22348	=>	60323,
		22349	=>	60321,
		22350	=>	60319,
		22351	=>	60318,
		22352	=>	60316,
		22353	=>	60314,
		22354	=>	60313,
		22355	=>	60311,
		22356	=>	60309,
		22357	=>	60307,
		22358	=>	60306,
		22359	=>	60304,
		22360	=>	60302,
		22361	=>	60301,
		22362	=>	60299,
		22363	=>	60297,
		22364	=>	60296,
		22365	=>	60294,
		22366	=>	60292,
		22367	=>	60290,
		22368	=>	60289,
		22369	=>	60287,
		22370	=>	60285,
		22371	=>	60284,
		22372	=>	60282,
		22373	=>	60280,
		22374	=>	60278,
		22375	=>	60277,
		22376	=>	60275,
		22377	=>	60273,
		22378	=>	60272,
		22379	=>	60270,
		22380	=>	60268,
		22381	=>	60267,
		22382	=>	60265,
		22383	=>	60263,
		22384	=>	60261,
		22385	=>	60260,
		22386	=>	60258,
		22387	=>	60256,
		22388	=>	60255,
		22389	=>	60253,
		22390	=>	60251,
		22391	=>	60249,
		22392	=>	60248,
		22393	=>	60246,
		22394	=>	60244,
		22395	=>	60243,
		22396	=>	60241,
		22397	=>	60239,
		22398	=>	60237,
		22399	=>	60236,
		22400	=>	60234,
		22401	=>	60232,
		22402	=>	60231,
		22403	=>	60229,
		22404	=>	60227,
		22405	=>	60225,
		22406	=>	60224,
		22407	=>	60222,
		22408	=>	60220,
		22409	=>	60219,
		22410	=>	60217,
		22411	=>	60215,
		22412	=>	60213,
		22413	=>	60212,
		22414	=>	60210,
		22415	=>	60208,
		22416	=>	60207,
		22417	=>	60205,
		22418	=>	60203,
		22419	=>	60201,
		22420	=>	60200,
		22421	=>	60198,
		22422	=>	60196,
		22423	=>	60195,
		22424	=>	60193,
		22425	=>	60191,
		22426	=>	60189,
		22427	=>	60188,
		22428	=>	60186,
		22429	=>	60184,
		22430	=>	60183,
		22431	=>	60181,
		22432	=>	60179,
		22433	=>	60177,
		22434	=>	60176,
		22435	=>	60174,
		22436	=>	60172,
		22437	=>	60170,
		22438	=>	60169,
		22439	=>	60167,
		22440	=>	60165,
		22441	=>	60164,
		22442	=>	60162,
		22443	=>	60160,
		22444	=>	60158,
		22445	=>	60157,
		22446	=>	60155,
		22447	=>	60153,
		22448	=>	60152,
		22449	=>	60150,
		22450	=>	60148,
		22451	=>	60146,
		22452	=>	60145,
		22453	=>	60143,
		22454	=>	60141,
		22455	=>	60139,
		22456	=>	60138,
		22457	=>	60136,
		22458	=>	60134,
		22459	=>	60133,
		22460	=>	60131,
		22461	=>	60129,
		22462	=>	60127,
		22463	=>	60126,
		22464	=>	60124,
		22465	=>	60122,
		22466	=>	60120,
		22467	=>	60119,
		22468	=>	60117,
		22469	=>	60115,
		22470	=>	60113,
		22471	=>	60112,
		22472	=>	60110,
		22473	=>	60108,
		22474	=>	60107,
		22475	=>	60105,
		22476	=>	60103,
		22477	=>	60101,
		22478	=>	60100,
		22479	=>	60098,
		22480	=>	60096,
		22481	=>	60094,
		22482	=>	60093,
		22483	=>	60091,
		22484	=>	60089,
		22485	=>	60087,
		22486	=>	60086,
		22487	=>	60084,
		22488	=>	60082,
		22489	=>	60081,
		22490	=>	60079,
		22491	=>	60077,
		22492	=>	60075,
		22493	=>	60074,
		22494	=>	60072,
		22495	=>	60070,
		22496	=>	60068,
		22497	=>	60067,
		22498	=>	60065,
		22499	=>	60063,
		22500	=>	60061,
		22501	=>	60060,
		22502	=>	60058,
		22503	=>	60056,
		22504	=>	60054,
		22505	=>	60053,
		22506	=>	60051,
		22507	=>	60049,
		22508	=>	60048,
		22509	=>	60046,
		22510	=>	60044,
		22511	=>	60042,
		22512	=>	60041,
		22513	=>	60039,
		22514	=>	60037,
		22515	=>	60035,
		22516	=>	60034,
		22517	=>	60032,
		22518	=>	60030,
		22519	=>	60028,
		22520	=>	60027,
		22521	=>	60025,
		22522	=>	60023,
		22523	=>	60021,
		22524	=>	60020,
		22525	=>	60018,
		22526	=>	60016,
		22527	=>	60014,
		22528	=>	60013,
		22529	=>	60011,
		22530	=>	60009,
		22531	=>	60007,
		22532	=>	60006,
		22533	=>	60004,
		22534	=>	60002,
		22535	=>	60000,
		22536	=>	59999,
		22537	=>	59997,
		22538	=>	59995,
		22539	=>	59993,
		22540	=>	59992,
		22541	=>	59990,
		22542	=>	59988,
		22543	=>	59986,
		22544	=>	59985,
		22545	=>	59983,
		22546	=>	59981,
		22547	=>	59979,
		22548	=>	59978,
		22549	=>	59976,
		22550	=>	59974,
		22551	=>	59972,
		22552	=>	59971,
		22553	=>	59969,
		22554	=>	59967,
		22555	=>	59965,
		22556	=>	59964,
		22557	=>	59962,
		22558	=>	59960,
		22559	=>	59958,
		22560	=>	59957,
		22561	=>	59955,
		22562	=>	59953,
		22563	=>	59951,
		22564	=>	59950,
		22565	=>	59948,
		22566	=>	59946,
		22567	=>	59944,
		22568	=>	59943,
		22569	=>	59941,
		22570	=>	59939,
		22571	=>	59937,
		22572	=>	59936,
		22573	=>	59934,
		22574	=>	59932,
		22575	=>	59930,
		22576	=>	59929,
		22577	=>	59927,
		22578	=>	59925,
		22579	=>	59923,
		22580	=>	59922,
		22581	=>	59920,
		22582	=>	59918,
		22583	=>	59916,
		22584	=>	59915,
		22585	=>	59913,
		22586	=>	59911,
		22587	=>	59909,
		22588	=>	59908,
		22589	=>	59906,
		22590	=>	59904,
		22591	=>	59902,
		22592	=>	59900,
		22593	=>	59899,
		22594	=>	59897,
		22595	=>	59895,
		22596	=>	59893,
		22597	=>	59892,
		22598	=>	59890,
		22599	=>	59888,
		22600	=>	59886,
		22601	=>	59885,
		22602	=>	59883,
		22603	=>	59881,
		22604	=>	59879,
		22605	=>	59878,
		22606	=>	59876,
		22607	=>	59874,
		22608	=>	59872,
		22609	=>	59870,
		22610	=>	59869,
		22611	=>	59867,
		22612	=>	59865,
		22613	=>	59863,
		22614	=>	59862,
		22615	=>	59860,
		22616	=>	59858,
		22617	=>	59856,
		22618	=>	59855,
		22619	=>	59853,
		22620	=>	59851,
		22621	=>	59849,
		22622	=>	59848,
		22623	=>	59846,
		22624	=>	59844,
		22625	=>	59842,
		22626	=>	59840,
		22627	=>	59839,
		22628	=>	59837,
		22629	=>	59835,
		22630	=>	59833,
		22631	=>	59832,
		22632	=>	59830,
		22633	=>	59828,
		22634	=>	59826,
		22635	=>	59824,
		22636	=>	59823,
		22637	=>	59821,
		22638	=>	59819,
		22639	=>	59817,
		22640	=>	59816,
		22641	=>	59814,
		22642	=>	59812,
		22643	=>	59810,
		22644	=>	59809,
		22645	=>	59807,
		22646	=>	59805,
		22647	=>	59803,
		22648	=>	59801,
		22649	=>	59800,
		22650	=>	59798,
		22651	=>	59796,
		22652	=>	59794,
		22653	=>	59793,
		22654	=>	59791,
		22655	=>	59789,
		22656	=>	59787,
		22657	=>	59785,
		22658	=>	59784,
		22659	=>	59782,
		22660	=>	59780,
		22661	=>	59778,
		22662	=>	59777,
		22663	=>	59775,
		22664	=>	59773,
		22665	=>	59771,
		22666	=>	59769,
		22667	=>	59768,
		22668	=>	59766,
		22669	=>	59764,
		22670	=>	59762,
		22671	=>	59761,
		22672	=>	59759,
		22673	=>	59757,
		22674	=>	59755,
		22675	=>	59753,
		22676	=>	59752,
		22677	=>	59750,
		22678	=>	59748,
		22679	=>	59746,
		22680	=>	59745,
		22681	=>	59743,
		22682	=>	59741,
		22683	=>	59739,
		22684	=>	59737,
		22685	=>	59736,
		22686	=>	59734,
		22687	=>	59732,
		22688	=>	59730,
		22689	=>	59728,
		22690	=>	59727,
		22691	=>	59725,
		22692	=>	59723,
		22693	=>	59721,
		22694	=>	59720,
		22695	=>	59718,
		22696	=>	59716,
		22697	=>	59714,
		22698	=>	59712,
		22699	=>	59711,
		22700	=>	59709,
		22701	=>	59707,
		22702	=>	59705,
		22703	=>	59703,
		22704	=>	59702,
		22705	=>	59700,
		22706	=>	59698,
		22707	=>	59696,
		22708	=>	59694,
		22709	=>	59693,
		22710	=>	59691,
		22711	=>	59689,
		22712	=>	59687,
		22713	=>	59686,
		22714	=>	59684,
		22715	=>	59682,
		22716	=>	59680,
		22717	=>	59678,
		22718	=>	59677,
		22719	=>	59675,
		22720	=>	59673,
		22721	=>	59671,
		22722	=>	59669,
		22723	=>	59668,
		22724	=>	59666,
		22725	=>	59664,
		22726	=>	59662,
		22727	=>	59660,
		22728	=>	59659,
		22729	=>	59657,
		22730	=>	59655,
		22731	=>	59653,
		22732	=>	59651,
		22733	=>	59650,
		22734	=>	59648,
		22735	=>	59646,
		22736	=>	59644,
		22737	=>	59642,
		22738	=>	59641,
		22739	=>	59639,
		22740	=>	59637,
		22741	=>	59635,
		22742	=>	59633,
		22743	=>	59632,
		22744	=>	59630,
		22745	=>	59628,
		22746	=>	59626,
		22747	=>	59624,
		22748	=>	59623,
		22749	=>	59621,
		22750	=>	59619,
		22751	=>	59617,
		22752	=>	59615,
		22753	=>	59614,
		22754	=>	59612,
		22755	=>	59610,
		22756	=>	59608,
		22757	=>	59606,
		22758	=>	59605,
		22759	=>	59603,
		22760	=>	59601,
		22761	=>	59599,
		22762	=>	59597,
		22763	=>	59596,
		22764	=>	59594,
		22765	=>	59592,
		22766	=>	59590,
		22767	=>	59588,
		22768	=>	59587,
		22769	=>	59585,
		22770	=>	59583,
		22771	=>	59581,
		22772	=>	59579,
		22773	=>	59578,
		22774	=>	59576,
		22775	=>	59574,
		22776	=>	59572,
		22777	=>	59570,
		22778	=>	59569,
		22779	=>	59567,
		22780	=>	59565,
		22781	=>	59563,
		22782	=>	59561,
		22783	=>	59560,
		22784	=>	59558,
		22785	=>	59556,
		22786	=>	59554,
		22787	=>	59552,
		22788	=>	59550,
		22789	=>	59549,
		22790	=>	59547,
		22791	=>	59545,
		22792	=>	59543,
		22793	=>	59541,
		22794	=>	59540,
		22795	=>	59538,
		22796	=>	59536,
		22797	=>	59534,
		22798	=>	59532,
		22799	=>	59531,
		22800	=>	59529,
		22801	=>	59527,
		22802	=>	59525,
		22803	=>	59523,
		22804	=>	59521,
		22805	=>	59520,
		22806	=>	59518,
		22807	=>	59516,
		22808	=>	59514,
		22809	=>	59512,
		22810	=>	59511,
		22811	=>	59509,
		22812	=>	59507,
		22813	=>	59505,
		22814	=>	59503,
		22815	=>	59502,
		22816	=>	59500,
		22817	=>	59498,
		22818	=>	59496,
		22819	=>	59494,
		22820	=>	59492,
		22821	=>	59491,
		22822	=>	59489,
		22823	=>	59487,
		22824	=>	59485,
		22825	=>	59483,
		22826	=>	59482,
		22827	=>	59480,
		22828	=>	59478,
		22829	=>	59476,
		22830	=>	59474,
		22831	=>	59472,
		22832	=>	59471,
		22833	=>	59469,
		22834	=>	59467,
		22835	=>	59465,
		22836	=>	59463,
		22837	=>	59461,
		22838	=>	59460,
		22839	=>	59458,
		22840	=>	59456,
		22841	=>	59454,
		22842	=>	59452,
		22843	=>	59451,
		22844	=>	59449,
		22845	=>	59447,
		22846	=>	59445,
		22847	=>	59443,
		22848	=>	59441,
		22849	=>	59440,
		22850	=>	59438,
		22851	=>	59436,
		22852	=>	59434,
		22853	=>	59432,
		22854	=>	59430,
		22855	=>	59429,
		22856	=>	59427,
		22857	=>	59425,
		22858	=>	59423,
		22859	=>	59421,
		22860	=>	59420,
		22861	=>	59418,
		22862	=>	59416,
		22863	=>	59414,
		22864	=>	59412,
		22865	=>	59410,
		22866	=>	59409,
		22867	=>	59407,
		22868	=>	59405,
		22869	=>	59403,
		22870	=>	59401,
		22871	=>	59399,
		22872	=>	59398,
		22873	=>	59396,
		22874	=>	59394,
		22875	=>	59392,
		22876	=>	59390,
		22877	=>	59388,
		22878	=>	59387,
		22879	=>	59385,
		22880	=>	59383,
		22881	=>	59381,
		22882	=>	59379,
		22883	=>	59377,
		22884	=>	59376,
		22885	=>	59374,
		22886	=>	59372,
		22887	=>	59370,
		22888	=>	59368,
		22889	=>	59366,
		22890	=>	59365,
		22891	=>	59363,
		22892	=>	59361,
		22893	=>	59359,
		22894	=>	59357,
		22895	=>	59355,
		22896	=>	59354,
		22897	=>	59352,
		22898	=>	59350,
		22899	=>	59348,
		22900	=>	59346,
		22901	=>	59344,
		22902	=>	59343,
		22903	=>	59341,
		22904	=>	59339,
		22905	=>	59337,
		22906	=>	59335,
		22907	=>	59333,
		22908	=>	59332,
		22909	=>	59330,
		22910	=>	59328,
		22911	=>	59326,
		22912	=>	59324,
		22913	=>	59322,
		22914	=>	59320,
		22915	=>	59319,
		22916	=>	59317,
		22917	=>	59315,
		22918	=>	59313,
		22919	=>	59311,
		22920	=>	59309,
		22921	=>	59308,
		22922	=>	59306,
		22923	=>	59304,
		22924	=>	59302,
		22925	=>	59300,
		22926	=>	59298,
		22927	=>	59297,
		22928	=>	59295,
		22929	=>	59293,
		22930	=>	59291,
		22931	=>	59289,
		22932	=>	59287,
		22933	=>	59285,
		22934	=>	59284,
		22935	=>	59282,
		22936	=>	59280,
		22937	=>	59278,
		22938	=>	59276,
		22939	=>	59274,
		22940	=>	59273,
		22941	=>	59271,
		22942	=>	59269,
		22943	=>	59267,
		22944	=>	59265,
		22945	=>	59263,
		22946	=>	59261,
		22947	=>	59260,
		22948	=>	59258,
		22949	=>	59256,
		22950	=>	59254,
		22951	=>	59252,
		22952	=>	59250,
		22953	=>	59248,
		22954	=>	59247,
		22955	=>	59245,
		22956	=>	59243,
		22957	=>	59241,
		22958	=>	59239,
		22959	=>	59237,
		22960	=>	59236,
		22961	=>	59234,
		22962	=>	59232,
		22963	=>	59230,
		22964	=>	59228,
		22965	=>	59226,
		22966	=>	59224,
		22967	=>	59223,
		22968	=>	59221,
		22969	=>	59219,
		22970	=>	59217,
		22971	=>	59215,
		22972	=>	59213,
		22973	=>	59211,
		22974	=>	59210,
		22975	=>	59208,
		22976	=>	59206,
		22977	=>	59204,
		22978	=>	59202,
		22979	=>	59200,
		22980	=>	59198,
		22981	=>	59197,
		22982	=>	59195,
		22983	=>	59193,
		22984	=>	59191,
		22985	=>	59189,
		22986	=>	59187,
		22987	=>	59185,
		22988	=>	59184,
		22989	=>	59182,
		22990	=>	59180,
		22991	=>	59178,
		22992	=>	59176,
		22993	=>	59174,
		22994	=>	59172,
		22995	=>	59171,
		22996	=>	59169,
		22997	=>	59167,
		22998	=>	59165,
		22999	=>	59163,
		23000	=>	59161,
		23001	=>	59159,
		23002	=>	59158,
		23003	=>	59156,
		23004	=>	59154,
		23005	=>	59152,
		23006	=>	59150,
		23007	=>	59148,
		23008	=>	59146,
		23009	=>	59145,
		23010	=>	59143,
		23011	=>	59141,
		23012	=>	59139,
		23013	=>	59137,
		23014	=>	59135,
		23015	=>	59133,
		23016	=>	59131,
		23017	=>	59130,
		23018	=>	59128,
		23019	=>	59126,
		23020	=>	59124,
		23021	=>	59122,
		23022	=>	59120,
		23023	=>	59118,
		23024	=>	59117,
		23025	=>	59115,
		23026	=>	59113,
		23027	=>	59111,
		23028	=>	59109,
		23029	=>	59107,
		23030	=>	59105,
		23031	=>	59103,
		23032	=>	59102,
		23033	=>	59100,
		23034	=>	59098,
		23035	=>	59096,
		23036	=>	59094,
		23037	=>	59092,
		23038	=>	59090,
		23039	=>	59088,
		23040	=>	59087,
		23041	=>	59085,
		23042	=>	59083,
		23043	=>	59081,
		23044	=>	59079,
		23045	=>	59077,
		23046	=>	59075,
		23047	=>	59073,
		23048	=>	59072,
		23049	=>	59070,
		23050	=>	59068,
		23051	=>	59066,
		23052	=>	59064,
		23053	=>	59062,
		23054	=>	59060,
		23055	=>	59059,
		23056	=>	59057,
		23057	=>	59055,
		23058	=>	59053,
		23059	=>	59051,
		23060	=>	59049,
		23061	=>	59047,
		23062	=>	59045,
		23063	=>	59043,
		23064	=>	59042,
		23065	=>	59040,
		23066	=>	59038,
		23067	=>	59036,
		23068	=>	59034,
		23069	=>	59032,
		23070	=>	59030,
		23071	=>	59028,
		23072	=>	59027,
		23073	=>	59025,
		23074	=>	59023,
		23075	=>	59021,
		23076	=>	59019,
		23077	=>	59017,
		23078	=>	59015,
		23079	=>	59013,
		23080	=>	59012,
		23081	=>	59010,
		23082	=>	59008,
		23083	=>	59006,
		23084	=>	59004,
		23085	=>	59002,
		23086	=>	59000,
		23087	=>	58998,
		23088	=>	58996,
		23089	=>	58995,
		23090	=>	58993,
		23091	=>	58991,
		23092	=>	58989,
		23093	=>	58987,
		23094	=>	58985,
		23095	=>	58983,
		23096	=>	58981,
		23097	=>	58980,
		23098	=>	58978,
		23099	=>	58976,
		23100	=>	58974,
		23101	=>	58972,
		23102	=>	58970,
		23103	=>	58968,
		23104	=>	58966,
		23105	=>	58964,
		23106	=>	58963,
		23107	=>	58961,
		23108	=>	58959,
		23109	=>	58957,
		23110	=>	58955,
		23111	=>	58953,
		23112	=>	58951,
		23113	=>	58949,
		23114	=>	58947,
		23115	=>	58946,
		23116	=>	58944,
		23117	=>	58942,
		23118	=>	58940,
		23119	=>	58938,
		23120	=>	58936,
		23121	=>	58934,
		23122	=>	58932,
		23123	=>	58930,
		23124	=>	58929,
		23125	=>	58927,
		23126	=>	58925,
		23127	=>	58923,
		23128	=>	58921,
		23129	=>	58919,
		23130	=>	58917,
		23131	=>	58915,
		23132	=>	58913,
		23133	=>	58912,
		23134	=>	58910,
		23135	=>	58908,
		23136	=>	58906,
		23137	=>	58904,
		23138	=>	58902,
		23139	=>	58900,
		23140	=>	58898,
		23141	=>	58896,
		23142	=>	58894,
		23143	=>	58893,
		23144	=>	58891,
		23145	=>	58889,
		23146	=>	58887,
		23147	=>	58885,
		23148	=>	58883,
		23149	=>	58881,
		23150	=>	58879,
		23151	=>	58877,
		23152	=>	58875,
		23153	=>	58874,
		23154	=>	58872,
		23155	=>	58870,
		23156	=>	58868,
		23157	=>	58866,
		23158	=>	58864,
		23159	=>	58862,
		23160	=>	58860,
		23161	=>	58858,
		23162	=>	58856,
		23163	=>	58855,
		23164	=>	58853,
		23165	=>	58851,
		23166	=>	58849,
		23167	=>	58847,
		23168	=>	58845,
		23169	=>	58843,
		23170	=>	58841,
		23171	=>	58839,
		23172	=>	58837,
		23173	=>	58836,
		23174	=>	58834,
		23175	=>	58832,
		23176	=>	58830,
		23177	=>	58828,
		23178	=>	58826,
		23179	=>	58824,
		23180	=>	58822,
		23181	=>	58820,
		23182	=>	58818,
		23183	=>	58817,
		23184	=>	58815,
		23185	=>	58813,
		23186	=>	58811,
		23187	=>	58809,
		23188	=>	58807,
		23189	=>	58805,
		23190	=>	58803,
		23191	=>	58801,
		23192	=>	58799,
		23193	=>	58797,
		23194	=>	58796,
		23195	=>	58794,
		23196	=>	58792,
		23197	=>	58790,
		23198	=>	58788,
		23199	=>	58786,
		23200	=>	58784,
		23201	=>	58782,
		23202	=>	58780,
		23203	=>	58778,
		23204	=>	58776,
		23205	=>	58775,
		23206	=>	58773,
		23207	=>	58771,
		23208	=>	58769,
		23209	=>	58767,
		23210	=>	58765,
		23211	=>	58763,
		23212	=>	58761,
		23213	=>	58759,
		23214	=>	58757,
		23215	=>	58755,
		23216	=>	58754,
		23217	=>	58752,
		23218	=>	58750,
		23219	=>	58748,
		23220	=>	58746,
		23221	=>	58744,
		23222	=>	58742,
		23223	=>	58740,
		23224	=>	58738,
		23225	=>	58736,
		23226	=>	58734,
		23227	=>	58732,
		23228	=>	58731,
		23229	=>	58729,
		23230	=>	58727,
		23231	=>	58725,
		23232	=>	58723,
		23233	=>	58721,
		23234	=>	58719,
		23235	=>	58717,
		23236	=>	58715,
		23237	=>	58713,
		23238	=>	58711,
		23239	=>	58709,
		23240	=>	58708,
		23241	=>	58706,
		23242	=>	58704,
		23243	=>	58702,
		23244	=>	58700,
		23245	=>	58698,
		23246	=>	58696,
		23247	=>	58694,
		23248	=>	58692,
		23249	=>	58690,
		23250	=>	58688,
		23251	=>	58686,
		23252	=>	58684,
		23253	=>	58683,
		23254	=>	58681,
		23255	=>	58679,
		23256	=>	58677,
		23257	=>	58675,
		23258	=>	58673,
		23259	=>	58671,
		23260	=>	58669,
		23261	=>	58667,
		23262	=>	58665,
		23263	=>	58663,
		23264	=>	58661,
		23265	=>	58659,
		23266	=>	58658,
		23267	=>	58656,
		23268	=>	58654,
		23269	=>	58652,
		23270	=>	58650,
		23271	=>	58648,
		23272	=>	58646,
		23273	=>	58644,
		23274	=>	58642,
		23275	=>	58640,
		23276	=>	58638,
		23277	=>	58636,
		23278	=>	58634,
		23279	=>	58632,
		23280	=>	58631,
		23281	=>	58629,
		23282	=>	58627,
		23283	=>	58625,
		23284	=>	58623,
		23285	=>	58621,
		23286	=>	58619,
		23287	=>	58617,
		23288	=>	58615,
		23289	=>	58613,
		23290	=>	58611,
		23291	=>	58609,
		23292	=>	58607,
		23293	=>	58605,
		23294	=>	58604,
		23295	=>	58602,
		23296	=>	58600,
		23297	=>	58598,
		23298	=>	58596,
		23299	=>	58594,
		23300	=>	58592,
		23301	=>	58590,
		23302	=>	58588,
		23303	=>	58586,
		23304	=>	58584,
		23305	=>	58582,
		23306	=>	58580,
		23307	=>	58578,
		23308	=>	58576,
		23309	=>	58574,
		23310	=>	58573,
		23311	=>	58571,
		23312	=>	58569,
		23313	=>	58567,
		23314	=>	58565,
		23315	=>	58563,
		23316	=>	58561,
		23317	=>	58559,
		23318	=>	58557,
		23319	=>	58555,
		23320	=>	58553,
		23321	=>	58551,
		23322	=>	58549,
		23323	=>	58547,
		23324	=>	58545,
		23325	=>	58543,
		23326	=>	58542,
		23327	=>	58540,
		23328	=>	58538,
		23329	=>	58536,
		23330	=>	58534,
		23331	=>	58532,
		23332	=>	58530,
		23333	=>	58528,
		23334	=>	58526,
		23335	=>	58524,
		23336	=>	58522,
		23337	=>	58520,
		23338	=>	58518,
		23339	=>	58516,
		23340	=>	58514,
		23341	=>	58512,
		23342	=>	58510,
		23343	=>	58509,
		23344	=>	58507,
		23345	=>	58505,
		23346	=>	58503,
		23347	=>	58501,
		23348	=>	58499,
		23349	=>	58497,
		23350	=>	58495,
		23351	=>	58493,
		23352	=>	58491,
		23353	=>	58489,
		23354	=>	58487,
		23355	=>	58485,
		23356	=>	58483,
		23357	=>	58481,
		23358	=>	58479,
		23359	=>	58477,
		23360	=>	58475,
		23361	=>	58474,
		23362	=>	58472,
		23363	=>	58470,
		23364	=>	58468,
		23365	=>	58466,
		23366	=>	58464,
		23367	=>	58462,
		23368	=>	58460,
		23369	=>	58458,
		23370	=>	58456,
		23371	=>	58454,
		23372	=>	58452,
		23373	=>	58450,
		23374	=>	58448,
		23375	=>	58446,
		23376	=>	58444,
		23377	=>	58442,
		23378	=>	58440,
		23379	=>	58438,
		23380	=>	58436,
		23381	=>	58434,
		23382	=>	58433,
		23383	=>	58431,
		23384	=>	58429,
		23385	=>	58427,
		23386	=>	58425,
		23387	=>	58423,
		23388	=>	58421,
		23389	=>	58419,
		23390	=>	58417,
		23391	=>	58415,
		23392	=>	58413,
		23393	=>	58411,
		23394	=>	58409,
		23395	=>	58407,
		23396	=>	58405,
		23397	=>	58403,
		23398	=>	58401,
		23399	=>	58399,
		23400	=>	58397,
		23401	=>	58395,
		23402	=>	58393,
		23403	=>	58391,
		23404	=>	58390,
		23405	=>	58388,
		23406	=>	58386,
		23407	=>	58384,
		23408	=>	58382,
		23409	=>	58380,
		23410	=>	58378,
		23411	=>	58376,
		23412	=>	58374,
		23413	=>	58372,
		23414	=>	58370,
		23415	=>	58368,
		23416	=>	58366,
		23417	=>	58364,
		23418	=>	58362,
		23419	=>	58360,
		23420	=>	58358,
		23421	=>	58356,
		23422	=>	58354,
		23423	=>	58352,
		23424	=>	58350,
		23425	=>	58348,
		23426	=>	58346,
		23427	=>	58344,
		23428	=>	58342,
		23429	=>	58340,
		23430	=>	58339,
		23431	=>	58337,
		23432	=>	58335,
		23433	=>	58333,
		23434	=>	58331,
		23435	=>	58329,
		23436	=>	58327,
		23437	=>	58325,
		23438	=>	58323,
		23439	=>	58321,
		23440	=>	58319,
		23441	=>	58317,
		23442	=>	58315,
		23443	=>	58313,
		23444	=>	58311,
		23445	=>	58309,
		23446	=>	58307,
		23447	=>	58305,
		23448	=>	58303,
		23449	=>	58301,
		23450	=>	58299,
		23451	=>	58297,
		23452	=>	58295,
		23453	=>	58293,
		23454	=>	58291,
		23455	=>	58289,
		23456	=>	58287,
		23457	=>	58285,
		23458	=>	58283,
		23459	=>	58281,
		23460	=>	58279,
		23461	=>	58278,
		23462	=>	58276,
		23463	=>	58274,
		23464	=>	58272,
		23465	=>	58270,
		23466	=>	58268,
		23467	=>	58266,
		23468	=>	58264,
		23469	=>	58262,
		23470	=>	58260,
		23471	=>	58258,
		23472	=>	58256,
		23473	=>	58254,
		23474	=>	58252,
		23475	=>	58250,
		23476	=>	58248,
		23477	=>	58246,
		23478	=>	58244,
		23479	=>	58242,
		23480	=>	58240,
		23481	=>	58238,
		23482	=>	58236,
		23483	=>	58234,
		23484	=>	58232,
		23485	=>	58230,
		23486	=>	58228,
		23487	=>	58226,
		23488	=>	58224,
		23489	=>	58222,
		23490	=>	58220,
		23491	=>	58218,
		23492	=>	58216,
		23493	=>	58214,
		23494	=>	58212,
		23495	=>	58210,
		23496	=>	58208,
		23497	=>	58206,
		23498	=>	58204,
		23499	=>	58202,
		23500	=>	58200,
		23501	=>	58198,
		23502	=>	58196,
		23503	=>	58194,
		23504	=>	58193,
		23505	=>	58191,
		23506	=>	58189,
		23507	=>	58187,
		23508	=>	58185,
		23509	=>	58183,
		23510	=>	58181,
		23511	=>	58179,
		23512	=>	58177,
		23513	=>	58175,
		23514	=>	58173,
		23515	=>	58171,
		23516	=>	58169,
		23517	=>	58167,
		23518	=>	58165,
		23519	=>	58163,
		23520	=>	58161,
		23521	=>	58159,
		23522	=>	58157,
		23523	=>	58155,
		23524	=>	58153,
		23525	=>	58151,
		23526	=>	58149,
		23527	=>	58147,
		23528	=>	58145,
		23529	=>	58143,
		23530	=>	58141,
		23531	=>	58139,
		23532	=>	58137,
		23533	=>	58135,
		23534	=>	58133,
		23535	=>	58131,
		23536	=>	58129,
		23537	=>	58127,
		23538	=>	58125,
		23539	=>	58123,
		23540	=>	58121,
		23541	=>	58119,
		23542	=>	58117,
		23543	=>	58115,
		23544	=>	58113,
		23545	=>	58111,
		23546	=>	58109,
		23547	=>	58107,
		23548	=>	58105,
		23549	=>	58103,
		23550	=>	58101,
		23551	=>	58099,
		23552	=>	58097,
		23553	=>	58095,
		23554	=>	58093,
		23555	=>	58091,
		23556	=>	58089,
		23557	=>	58087,
		23558	=>	58085,
		23559	=>	58083,
		23560	=>	58081,
		23561	=>	58079,
		23562	=>	58077,
		23563	=>	58075,
		23564	=>	58073,
		23565	=>	58071,
		23566	=>	58069,
		23567	=>	58067,
		23568	=>	58065,
		23569	=>	58063,
		23570	=>	58061,
		23571	=>	58059,
		23572	=>	58057,
		23573	=>	58055,
		23574	=>	58053,
		23575	=>	58051,
		23576	=>	58049,
		23577	=>	58047,
		23578	=>	58045,
		23579	=>	58043,
		23580	=>	58041,
		23581	=>	58039,
		23582	=>	58037,
		23583	=>	58035,
		23584	=>	58033,
		23585	=>	58031,
		23586	=>	58029,
		23587	=>	58027,
		23588	=>	58025,
		23589	=>	58023,
		23590	=>	58021,
		23591	=>	58019,
		23592	=>	58017,
		23593	=>	58015,
		23594	=>	58013,
		23595	=>	58011,
		23596	=>	58009,
		23597	=>	58007,
		23598	=>	58005,
		23599	=>	58003,
		23600	=>	58001,
		23601	=>	57999,
		23602	=>	57997,
		23603	=>	57995,
		23604	=>	57993,
		23605	=>	57991,
		23606	=>	57989,
		23607	=>	57987,
		23608	=>	57985,
		23609	=>	57983,
		23610	=>	57981,
		23611	=>	57979,
		23612	=>	57977,
		23613	=>	57975,
		23614	=>	57973,
		23615	=>	57971,
		23616	=>	57969,
		23617	=>	57967,
		23618	=>	57965,
		23619	=>	57963,
		23620	=>	57961,
		23621	=>	57959,
		23622	=>	57957,
		23623	=>	57955,
		23624	=>	57953,
		23625	=>	57951,
		23626	=>	57949,
		23627	=>	57947,
		23628	=>	57945,
		23629	=>	57943,
		23630	=>	57941,
		23631	=>	57939,
		23632	=>	57937,
		23633	=>	57935,
		23634	=>	57933,
		23635	=>	57931,
		23636	=>	57929,
		23637	=>	57927,
		23638	=>	57925,
		23639	=>	57923,
		23640	=>	57921,
		23641	=>	57919,
		23642	=>	57917,
		23643	=>	57915,
		23644	=>	57913,
		23645	=>	57911,
		23646	=>	57909,
		23647	=>	57907,
		23648	=>	57905,
		23649	=>	57903,
		23650	=>	57901,
		23651	=>	57899,
		23652	=>	57897,
		23653	=>	57895,
		23654	=>	57893,
		23655	=>	57891,
		23656	=>	57889,
		23657	=>	57887,
		23658	=>	57885,
		23659	=>	57883,
		23660	=>	57881,
		23661	=>	57879,
		23662	=>	57876,
		23663	=>	57874,
		23664	=>	57872,
		23665	=>	57870,
		23666	=>	57868,
		23667	=>	57866,
		23668	=>	57864,
		23669	=>	57862,
		23670	=>	57860,
		23671	=>	57858,
		23672	=>	57856,
		23673	=>	57854,
		23674	=>	57852,
		23675	=>	57850,
		23676	=>	57848,
		23677	=>	57846,
		23678	=>	57844,
		23679	=>	57842,
		23680	=>	57840,
		23681	=>	57838,
		23682	=>	57836,
		23683	=>	57834,
		23684	=>	57832,
		23685	=>	57830,
		23686	=>	57828,
		23687	=>	57826,
		23688	=>	57824,
		23689	=>	57822,
		23690	=>	57820,
		23691	=>	57818,
		23692	=>	57816,
		23693	=>	57814,
		23694	=>	57812,
		23695	=>	57810,
		23696	=>	57808,
		23697	=>	57806,
		23698	=>	57804,
		23699	=>	57802,
		23700	=>	57800,
		23701	=>	57798,
		23702	=>	57796,
		23703	=>	57794,
		23704	=>	57792,
		23705	=>	57789,
		23706	=>	57787,
		23707	=>	57785,
		23708	=>	57783,
		23709	=>	57781,
		23710	=>	57779,
		23711	=>	57777,
		23712	=>	57775,
		23713	=>	57773,
		23714	=>	57771,
		23715	=>	57769,
		23716	=>	57767,
		23717	=>	57765,
		23718	=>	57763,
		23719	=>	57761,
		23720	=>	57759,
		23721	=>	57757,
		23722	=>	57755,
		23723	=>	57753,
		23724	=>	57751,
		23725	=>	57749,
		23726	=>	57747,
		23727	=>	57745,
		23728	=>	57743,
		23729	=>	57741,
		23730	=>	57739,
		23731	=>	57737,
		23732	=>	57735,
		23733	=>	57733,
		23734	=>	57731,
		23735	=>	57729,
		23736	=>	57726,
		23737	=>	57724,
		23738	=>	57722,
		23739	=>	57720,
		23740	=>	57718,
		23741	=>	57716,
		23742	=>	57714,
		23743	=>	57712,
		23744	=>	57710,
		23745	=>	57708,
		23746	=>	57706,
		23747	=>	57704,
		23748	=>	57702,
		23749	=>	57700,
		23750	=>	57698,
		23751	=>	57696,
		23752	=>	57694,
		23753	=>	57692,
		23754	=>	57690,
		23755	=>	57688,
		23756	=>	57686,
		23757	=>	57684,
		23758	=>	57682,
		23759	=>	57680,
		23760	=>	57678,
		23761	=>	57676,
		23762	=>	57673,
		23763	=>	57671,
		23764	=>	57669,
		23765	=>	57667,
		23766	=>	57665,
		23767	=>	57663,
		23768	=>	57661,
		23769	=>	57659,
		23770	=>	57657,
		23771	=>	57655,
		23772	=>	57653,
		23773	=>	57651,
		23774	=>	57649,
		23775	=>	57647,
		23776	=>	57645,
		23777	=>	57643,
		23778	=>	57641,
		23779	=>	57639,
		23780	=>	57637,
		23781	=>	57635,
		23782	=>	57633,
		23783	=>	57631,
		23784	=>	57629,
		23785	=>	57626,
		23786	=>	57624,
		23787	=>	57622,
		23788	=>	57620,
		23789	=>	57618,
		23790	=>	57616,
		23791	=>	57614,
		23792	=>	57612,
		23793	=>	57610,
		23794	=>	57608,
		23795	=>	57606,
		23796	=>	57604,
		23797	=>	57602,
		23798	=>	57600,
		23799	=>	57598,
		23800	=>	57596,
		23801	=>	57594,
		23802	=>	57592,
		23803	=>	57590,
		23804	=>	57588,
		23805	=>	57585,
		23806	=>	57583,
		23807	=>	57581,
		23808	=>	57579,
		23809	=>	57577,
		23810	=>	57575,
		23811	=>	57573,
		23812	=>	57571,
		23813	=>	57569,
		23814	=>	57567,
		23815	=>	57565,
		23816	=>	57563,
		23817	=>	57561,
		23818	=>	57559,
		23819	=>	57557,
		23820	=>	57555,
		23821	=>	57553,
		23822	=>	57551,
		23823	=>	57549,
		23824	=>	57546,
		23825	=>	57544,
		23826	=>	57542,
		23827	=>	57540,
		23828	=>	57538,
		23829	=>	57536,
		23830	=>	57534,
		23831	=>	57532,
		23832	=>	57530,
		23833	=>	57528,
		23834	=>	57526,
		23835	=>	57524,
		23836	=>	57522,
		23837	=>	57520,
		23838	=>	57518,
		23839	=>	57516,
		23840	=>	57514,
		23841	=>	57512,
		23842	=>	57509,
		23843	=>	57507,
		23844	=>	57505,
		23845	=>	57503,
		23846	=>	57501,
		23847	=>	57499,
		23848	=>	57497,
		23849	=>	57495,
		23850	=>	57493,
		23851	=>	57491,
		23852	=>	57489,
		23853	=>	57487,
		23854	=>	57485,
		23855	=>	57483,
		23856	=>	57481,
		23857	=>	57479,
		23858	=>	57476,
		23859	=>	57474,
		23860	=>	57472,
		23861	=>	57470,
		23862	=>	57468,
		23863	=>	57466,
		23864	=>	57464,
		23865	=>	57462,
		23866	=>	57460,
		23867	=>	57458,
		23868	=>	57456,
		23869	=>	57454,
		23870	=>	57452,
		23871	=>	57450,
		23872	=>	57448,
		23873	=>	57445,
		23874	=>	57443,
		23875	=>	57441,
		23876	=>	57439,
		23877	=>	57437,
		23878	=>	57435,
		23879	=>	57433,
		23880	=>	57431,
		23881	=>	57429,
		23882	=>	57427,
		23883	=>	57425,
		23884	=>	57423,
		23885	=>	57421,
		23886	=>	57419,
		23887	=>	57417,
		23888	=>	57414,
		23889	=>	57412,
		23890	=>	57410,
		23891	=>	57408,
		23892	=>	57406,
		23893	=>	57404,
		23894	=>	57402,
		23895	=>	57400,
		23896	=>	57398,
		23897	=>	57396,
		23898	=>	57394,
		23899	=>	57392,
		23900	=>	57390,
		23901	=>	57388,
		23902	=>	57385,
		23903	=>	57383,
		23904	=>	57381,
		23905	=>	57379,
		23906	=>	57377,
		23907	=>	57375,
		23908	=>	57373,
		23909	=>	57371,
		23910	=>	57369,
		23911	=>	57367,
		23912	=>	57365,
		23913	=>	57363,
		23914	=>	57361,
		23915	=>	57358,
		23916	=>	57356,
		23917	=>	57354,
		23918	=>	57352,
		23919	=>	57350,
		23920	=>	57348,
		23921	=>	57346,
		23922	=>	57344,
		23923	=>	57342,
		23924	=>	57340,
		23925	=>	57338,
		23926	=>	57336,
		23927	=>	57334,
		23928	=>	57331,
		23929	=>	57329,
		23930	=>	57327,
		23931	=>	57325,
		23932	=>	57323,
		23933	=>	57321,
		23934	=>	57319,
		23935	=>	57317,
		23936	=>	57315,
		23937	=>	57313,
		23938	=>	57311,
		23939	=>	57309,
		23940	=>	57307,
		23941	=>	57304,
		23942	=>	57302,
		23943	=>	57300,
		23944	=>	57298,
		23945	=>	57296,
		23946	=>	57294,
		23947	=>	57292,
		23948	=>	57290,
		23949	=>	57288,
		23950	=>	57286,
		23951	=>	57284,
		23952	=>	57282,
		23953	=>	57279,
		23954	=>	57277,
		23955	=>	57275,
		23956	=>	57273,
		23957	=>	57271,
		23958	=>	57269,
		23959	=>	57267,
		23960	=>	57265,
		23961	=>	57263,
		23962	=>	57261,
		23963	=>	57259,
		23964	=>	57256,
		23965	=>	57254,
		23966	=>	57252,
		23967	=>	57250,
		23968	=>	57248,
		23969	=>	57246,
		23970	=>	57244,
		23971	=>	57242,
		23972	=>	57240,
		23973	=>	57238,
		23974	=>	57236,
		23975	=>	57233,
		23976	=>	57231,
		23977	=>	57229,
		23978	=>	57227,
		23979	=>	57225,
		23980	=>	57223,
		23981	=>	57221,
		23982	=>	57219,
		23983	=>	57217,
		23984	=>	57215,
		23985	=>	57213,
		23986	=>	57210,
		23987	=>	57208,
		23988	=>	57206,
		23989	=>	57204,
		23990	=>	57202,
		23991	=>	57200,
		23992	=>	57198,
		23993	=>	57196,
		23994	=>	57194,
		23995	=>	57192,
		23996	=>	57190,
		23997	=>	57187,
		23998	=>	57185,
		23999	=>	57183,
		24000	=>	57181,
		24001	=>	57179,
		24002	=>	57177,
		24003	=>	57175,
		24004	=>	57173,
		24005	=>	57171,
		24006	=>	57169,
		24007	=>	57167,
		24008	=>	57164,
		24009	=>	57162,
		24010	=>	57160,
		24011	=>	57158,
		24012	=>	57156,
		24013	=>	57154,
		24014	=>	57152,
		24015	=>	57150,
		24016	=>	57148,
		24017	=>	57146,
		24018	=>	57143,
		24019	=>	57141,
		24020	=>	57139,
		24021	=>	57137,
		24022	=>	57135,
		24023	=>	57133,
		24024	=>	57131,
		24025	=>	57129,
		24026	=>	57127,
		24027	=>	57125,
		24028	=>	57122,
		24029	=>	57120,
		24030	=>	57118,
		24031	=>	57116,
		24032	=>	57114,
		24033	=>	57112,
		24034	=>	57110,
		24035	=>	57108,
		24036	=>	57106,
		24037	=>	57103,
		24038	=>	57101,
		24039	=>	57099,
		24040	=>	57097,
		24041	=>	57095,
		24042	=>	57093,
		24043	=>	57091,
		24044	=>	57089,
		24045	=>	57087,
		24046	=>	57085,
		24047	=>	57082,
		24048	=>	57080,
		24049	=>	57078,
		24050	=>	57076,
		24051	=>	57074,
		24052	=>	57072,
		24053	=>	57070,
		24054	=>	57068,
		24055	=>	57066,
		24056	=>	57063,
		24057	=>	57061,
		24058	=>	57059,
		24059	=>	57057,
		24060	=>	57055,
		24061	=>	57053,
		24062	=>	57051,
		24063	=>	57049,
		24064	=>	57047,
		24065	=>	57045,
		24066	=>	57042,
		24067	=>	57040,
		24068	=>	57038,
		24069	=>	57036,
		24070	=>	57034,
		24071	=>	57032,
		24072	=>	57030,
		24073	=>	57028,
		24074	=>	57026,
		24075	=>	57023,
		24076	=>	57021,
		24077	=>	57019,
		24078	=>	57017,
		24079	=>	57015,
		24080	=>	57013,
		24081	=>	57011,
		24082	=>	57009,
		24083	=>	57006,
		24084	=>	57004,
		24085	=>	57002,
		24086	=>	57000,
		24087	=>	56998,
		24088	=>	56996,
		24089	=>	56994,
		24090	=>	56992,
		24091	=>	56990,
		24092	=>	56987,
		24093	=>	56985,
		24094	=>	56983,
		24095	=>	56981,
		24096	=>	56979,
		24097	=>	56977,
		24098	=>	56975,
		24099	=>	56973,
		24100	=>	56971,
		24101	=>	56968,
		24102	=>	56966,
		24103	=>	56964,
		24104	=>	56962,
		24105	=>	56960,
		24106	=>	56958,
		24107	=>	56956,
		24108	=>	56954,
		24109	=>	56951,
		24110	=>	56949,
		24111	=>	56947,
		24112	=>	56945,
		24113	=>	56943,
		24114	=>	56941,
		24115	=>	56939,
		24116	=>	56937,
		24117	=>	56934,
		24118	=>	56932,
		24119	=>	56930,
		24120	=>	56928,
		24121	=>	56926,
		24122	=>	56924,
		24123	=>	56922,
		24124	=>	56920,
		24125	=>	56918,
		24126	=>	56915,
		24127	=>	56913,
		24128	=>	56911,
		24129	=>	56909,
		24130	=>	56907,
		24131	=>	56905,
		24132	=>	56903,
		24133	=>	56901,
		24134	=>	56898,
		24135	=>	56896,
		24136	=>	56894,
		24137	=>	56892,
		24138	=>	56890,
		24139	=>	56888,
		24140	=>	56886,
		24141	=>	56884,
		24142	=>	56881,
		24143	=>	56879,
		24144	=>	56877,
		24145	=>	56875,
		24146	=>	56873,
		24147	=>	56871,
		24148	=>	56869,
		24149	=>	56866,
		24150	=>	56864,
		24151	=>	56862,
		24152	=>	56860,
		24153	=>	56858,
		24154	=>	56856,
		24155	=>	56854,
		24156	=>	56852,
		24157	=>	56849,
		24158	=>	56847,
		24159	=>	56845,
		24160	=>	56843,
		24161	=>	56841,
		24162	=>	56839,
		24163	=>	56837,
		24164	=>	56835,
		24165	=>	56832,
		24166	=>	56830,
		24167	=>	56828,
		24168	=>	56826,
		24169	=>	56824,
		24170	=>	56822,
		24171	=>	56820,
		24172	=>	56817,
		24173	=>	56815,
		24174	=>	56813,
		24175	=>	56811,
		24176	=>	56809,
		24177	=>	56807,
		24178	=>	56805,
		24179	=>	56803,
		24180	=>	56800,
		24181	=>	56798,
		24182	=>	56796,
		24183	=>	56794,
		24184	=>	56792,
		24185	=>	56790,
		24186	=>	56788,
		24187	=>	56785,
		24188	=>	56783,
		24189	=>	56781,
		24190	=>	56779,
		24191	=>	56777,
		24192	=>	56775,
		24193	=>	56773,
		24194	=>	56770,
		24195	=>	56768,
		24196	=>	56766,
		24197	=>	56764,
		24198	=>	56762,
		24199	=>	56760,
		24200	=>	56758,
		24201	=>	56755,
		24202	=>	56753,
		24203	=>	56751,
		24204	=>	56749,
		24205	=>	56747,
		24206	=>	56745,
		24207	=>	56743,
		24208	=>	56741,
		24209	=>	56738,
		24210	=>	56736,
		24211	=>	56734,
		24212	=>	56732,
		24213	=>	56730,
		24214	=>	56728,
		24215	=>	56726,
		24216	=>	56723,
		24217	=>	56721,
		24218	=>	56719,
		24219	=>	56717,
		24220	=>	56715,
		24221	=>	56713,
		24222	=>	56711,
		24223	=>	56708,
		24224	=>	56706,
		24225	=>	56704,
		24226	=>	56702,
		24227	=>	56700,
		24228	=>	56698,
		24229	=>	56695,
		24230	=>	56693,
		24231	=>	56691,
		24232	=>	56689,
		24233	=>	56687,
		24234	=>	56685,
		24235	=>	56683,
		24236	=>	56680,
		24237	=>	56678,
		24238	=>	56676,
		24239	=>	56674,
		24240	=>	56672,
		24241	=>	56670,
		24242	=>	56668,
		24243	=>	56665,
		24244	=>	56663,
		24245	=>	56661,
		24246	=>	56659,
		24247	=>	56657,
		24248	=>	56655,
		24249	=>	56653,
		24250	=>	56650,
		24251	=>	56648,
		24252	=>	56646,
		24253	=>	56644,
		24254	=>	56642,
		24255	=>	56640,
		24256	=>	56637,
		24257	=>	56635,
		24258	=>	56633,
		24259	=>	56631,
		24260	=>	56629,
		24261	=>	56627,
		24262	=>	56625,
		24263	=>	56622,
		24264	=>	56620,
		24265	=>	56618,
		24266	=>	56616,
		24267	=>	56614,
		24268	=>	56612,
		24269	=>	56609,
		24270	=>	56607,
		24271	=>	56605,
		24272	=>	56603,
		24273	=>	56601,
		24274	=>	56599,
		24275	=>	56597,
		24276	=>	56594,
		24277	=>	56592,
		24278	=>	56590,
		24279	=>	56588,
		24280	=>	56586,
		24281	=>	56584,
		24282	=>	56581,
		24283	=>	56579,
		24284	=>	56577,
		24285	=>	56575,
		24286	=>	56573,
		24287	=>	56571,
		24288	=>	56568,
		24289	=>	56566,
		24290	=>	56564,
		24291	=>	56562,
		24292	=>	56560,
		24293	=>	56558,
		24294	=>	56556,
		24295	=>	56553,
		24296	=>	56551,
		24297	=>	56549,
		24298	=>	56547,
		24299	=>	56545,
		24300	=>	56543,
		24301	=>	56540,
		24302	=>	56538,
		24303	=>	56536,
		24304	=>	56534,
		24305	=>	56532,
		24306	=>	56530,
		24307	=>	56527,
		24308	=>	56525,
		24309	=>	56523,
		24310	=>	56521,
		24311	=>	56519,
		24312	=>	56517,
		24313	=>	56514,
		24314	=>	56512,
		24315	=>	56510,
		24316	=>	56508,
		24317	=>	56506,
		24318	=>	56504,
		24319	=>	56501,
		24320	=>	56499,
		24321	=>	56497,
		24322	=>	56495,
		24323	=>	56493,
		24324	=>	56491,
		24325	=>	56488,
		24326	=>	56486,
		24327	=>	56484,
		24328	=>	56482,
		24329	=>	56480,
		24330	=>	56478,
		24331	=>	56475,
		24332	=>	56473,
		24333	=>	56471,
		24334	=>	56469,
		24335	=>	56467,
		24336	=>	56465,
		24337	=>	56462,
		24338	=>	56460,
		24339	=>	56458,
		24340	=>	56456,
		24341	=>	56454,
		24342	=>	56452,
		24343	=>	56449,
		24344	=>	56447,
		24345	=>	56445,
		24346	=>	56443,
		24347	=>	56441,
		24348	=>	56439,
		24349	=>	56436,
		24350	=>	56434,
		24351	=>	56432,
		24352	=>	56430,
		24353	=>	56428,
		24354	=>	56425,
		24355	=>	56423,
		24356	=>	56421,
		24357	=>	56419,
		24358	=>	56417,
		24359	=>	56415,
		24360	=>	56412,
		24361	=>	56410,
		24362	=>	56408,
		24363	=>	56406,
		24364	=>	56404,
		24365	=>	56402,
		24366	=>	56399,
		24367	=>	56397,
		24368	=>	56395,
		24369	=>	56393,
		24370	=>	56391,
		24371	=>	56389,
		24372	=>	56386,
		24373	=>	56384,
		24374	=>	56382,
		24375	=>	56380,
		24376	=>	56378,
		24377	=>	56375,
		24378	=>	56373,
		24379	=>	56371,
		24380	=>	56369,
		24381	=>	56367,
		24382	=>	56365,
		24383	=>	56362,
		24384	=>	56360,
		24385	=>	56358,
		24386	=>	56356,
		24387	=>	56354,
		24388	=>	56351,
		24389	=>	56349,
		24390	=>	56347,
		24391	=>	56345,
		24392	=>	56343,
		24393	=>	56341,
		24394	=>	56338,
		24395	=>	56336,
		24396	=>	56334,
		24397	=>	56332,
		24398	=>	56330,
		24399	=>	56327,
		24400	=>	56325,
		24401	=>	56323,
		24402	=>	56321,
		24403	=>	56319,
		24404	=>	56317,
		24405	=>	56314,
		24406	=>	56312,
		24407	=>	56310,
		24408	=>	56308,
		24409	=>	56306,
		24410	=>	56303,
		24411	=>	56301,
		24412	=>	56299,
		24413	=>	56297,
		24414	=>	56295,
		24415	=>	56292,
		24416	=>	56290,
		24417	=>	56288,
		24418	=>	56286,
		24419	=>	56284,
		24420	=>	56282,
		24421	=>	56279,
		24422	=>	56277,
		24423	=>	56275,
		24424	=>	56273,
		24425	=>	56271,
		24426	=>	56268,
		24427	=>	56266,
		24428	=>	56264,
		24429	=>	56262,
		24430	=>	56260,
		24431	=>	56257,
		24432	=>	56255,
		24433	=>	56253,
		24434	=>	56251,
		24435	=>	56249,
		24436	=>	56247,
		24437	=>	56244,
		24438	=>	56242,
		24439	=>	56240,
		24440	=>	56238,
		24441	=>	56236,
		24442	=>	56233,
		24443	=>	56231,
		24444	=>	56229,
		24445	=>	56227,
		24446	=>	56225,
		24447	=>	56222,
		24448	=>	56220,
		24449	=>	56218,
		24450	=>	56216,
		24451	=>	56214,
		24452	=>	56211,
		24453	=>	56209,
		24454	=>	56207,
		24455	=>	56205,
		24456	=>	56203,
		24457	=>	56200,
		24458	=>	56198,
		24459	=>	56196,
		24460	=>	56194,
		24461	=>	56192,
		24462	=>	56189,
		24463	=>	56187,
		24464	=>	56185,
		24465	=>	56183,
		24466	=>	56181,
		24467	=>	56178,
		24468	=>	56176,
		24469	=>	56174,
		24470	=>	56172,
		24471	=>	56170,
		24472	=>	56167,
		24473	=>	56165,
		24474	=>	56163,
		24475	=>	56161,
		24476	=>	56159,
		24477	=>	56156,
		24478	=>	56154,
		24479	=>	56152,
		24480	=>	56150,
		24481	=>	56148,
		24482	=>	56145,
		24483	=>	56143,
		24484	=>	56141,
		24485	=>	56139,
		24486	=>	56137,
		24487	=>	56134,
		24488	=>	56132,
		24489	=>	56130,
		24490	=>	56128,
		24491	=>	56126,
		24492	=>	56123,
		24493	=>	56121,
		24494	=>	56119,
		24495	=>	56117,
		24496	=>	56115,
		24497	=>	56112,
		24498	=>	56110,
		24499	=>	56108,
		24500	=>	56106,
		24501	=>	56104,
		24502	=>	56101,
		24503	=>	56099,
		24504	=>	56097,
		24505	=>	56095,
		24506	=>	56093,
		24507	=>	56090,
		24508	=>	56088,
		24509	=>	56086,
		24510	=>	56084,
		24511	=>	56082,
		24512	=>	56079,
		24513	=>	56077,
		24514	=>	56075,
		24515	=>	56073,
		24516	=>	56071,
		24517	=>	56068,
		24518	=>	56066,
		24519	=>	56064,
		24520	=>	56062,
		24521	=>	56059,
		24522	=>	56057,
		24523	=>	56055,
		24524	=>	56053,
		24525	=>	56051,
		24526	=>	56048,
		24527	=>	56046,
		24528	=>	56044,
		24529	=>	56042,
		24530	=>	56040,
		24531	=>	56037,
		24532	=>	56035,
		24533	=>	56033,
		24534	=>	56031,
		24535	=>	56029,
		24536	=>	56026,
		24537	=>	56024,
		24538	=>	56022,
		24539	=>	56020,
		24540	=>	56017,
		24541	=>	56015,
		24542	=>	56013,
		24543	=>	56011,
		24544	=>	56009,
		24545	=>	56006,
		24546	=>	56004,
		24547	=>	56002,
		24548	=>	56000,
		24549	=>	55998,
		24550	=>	55995,
		24551	=>	55993,
		24552	=>	55991,
		24553	=>	55989,
		24554	=>	55986,
		24555	=>	55984,
		24556	=>	55982,
		24557	=>	55980,
		24558	=>	55978,
		24559	=>	55975,
		24560	=>	55973,
		24561	=>	55971,
		24562	=>	55969,
		24563	=>	55966,
		24564	=>	55964,
		24565	=>	55962,
		24566	=>	55960,
		24567	=>	55958,
		24568	=>	55955,
		24569	=>	55953,
		24570	=>	55951,
		24571	=>	55949,
		24572	=>	55947,
		24573	=>	55944,
		24574	=>	55942,
		24575	=>	55940,
		24576	=>	55938,
		24577	=>	55935,
		24578	=>	55933,
		24579	=>	55931,
		24580	=>	55929,
		24581	=>	55927,
		24582	=>	55924,
		24583	=>	55922,
		24584	=>	55920,
		24585	=>	55918,
		24586	=>	55915,
		24587	=>	55913,
		24588	=>	55911,
		24589	=>	55909,
		24590	=>	55907,
		24591	=>	55904,
		24592	=>	55902,
		24593	=>	55900,
		24594	=>	55898,
		24595	=>	55895,
		24596	=>	55893,
		24597	=>	55891,
		24598	=>	55889,
		24599	=>	55886,
		24600	=>	55884,
		24601	=>	55882,
		24602	=>	55880,
		24603	=>	55878,
		24604	=>	55875,
		24605	=>	55873,
		24606	=>	55871,
		24607	=>	55869,
		24608	=>	55866,
		24609	=>	55864,
		24610	=>	55862,
		24611	=>	55860,
		24612	=>	55858,
		24613	=>	55855,
		24614	=>	55853,
		24615	=>	55851,
		24616	=>	55849,
		24617	=>	55846,
		24618	=>	55844,
		24619	=>	55842,
		24620	=>	55840,
		24621	=>	55837,
		24622	=>	55835,
		24623	=>	55833,
		24624	=>	55831,
		24625	=>	55829,
		24626	=>	55826,
		24627	=>	55824,
		24628	=>	55822,
		24629	=>	55820,
		24630	=>	55817,
		24631	=>	55815,
		24632	=>	55813,
		24633	=>	55811,
		24634	=>	55808,
		24635	=>	55806,
		24636	=>	55804,
		24637	=>	55802,
		24638	=>	55799,
		24639	=>	55797,
		24640	=>	55795,
		24641	=>	55793,
		24642	=>	55791,
		24643	=>	55788,
		24644	=>	55786,
		24645	=>	55784,
		24646	=>	55782,
		24647	=>	55779,
		24648	=>	55777,
		24649	=>	55775,
		24650	=>	55773,
		24651	=>	55770,
		24652	=>	55768,
		24653	=>	55766,
		24654	=>	55764,
		24655	=>	55761,
		24656	=>	55759,
		24657	=>	55757,
		24658	=>	55755,
		24659	=>	55753,
		24660	=>	55750,
		24661	=>	55748,
		24662	=>	55746,
		24663	=>	55744,
		24664	=>	55741,
		24665	=>	55739,
		24666	=>	55737,
		24667	=>	55735,
		24668	=>	55732,
		24669	=>	55730,
		24670	=>	55728,
		24671	=>	55726,
		24672	=>	55723,
		24673	=>	55721,
		24674	=>	55719,
		24675	=>	55717,
		24676	=>	55714,
		24677	=>	55712,
		24678	=>	55710,
		24679	=>	55708,
		24680	=>	55705,
		24681	=>	55703,
		24682	=>	55701,
		24683	=>	55699,
		24684	=>	55696,
		24685	=>	55694,
		24686	=>	55692,
		24687	=>	55690,
		24688	=>	55687,
		24689	=>	55685,
		24690	=>	55683,
		24691	=>	55681,
		24692	=>	55679,
		24693	=>	55676,
		24694	=>	55674,
		24695	=>	55672,
		24696	=>	55670,
		24697	=>	55667,
		24698	=>	55665,
		24699	=>	55663,
		24700	=>	55661,
		24701	=>	55658,
		24702	=>	55656,
		24703	=>	55654,
		24704	=>	55652,
		24705	=>	55649,
		24706	=>	55647,
		24707	=>	55645,
		24708	=>	55643,
		24709	=>	55640,
		24710	=>	55638,
		24711	=>	55636,
		24712	=>	55634,
		24713	=>	55631,
		24714	=>	55629,
		24715	=>	55627,
		24716	=>	55625,
		24717	=>	55622,
		24718	=>	55620,
		24719	=>	55618,
		24720	=>	55616,
		24721	=>	55613,
		24722	=>	55611,
		24723	=>	55609,
		24724	=>	55607,
		24725	=>	55604,
		24726	=>	55602,
		24727	=>	55600,
		24728	=>	55598,
		24729	=>	55595,
		24730	=>	55593,
		24731	=>	55591,
		24732	=>	55589,
		24733	=>	55586,
		24734	=>	55584,
		24735	=>	55582,
		24736	=>	55579,
		24737	=>	55577,
		24738	=>	55575,
		24739	=>	55573,
		24740	=>	55570,
		24741	=>	55568,
		24742	=>	55566,
		24743	=>	55564,
		24744	=>	55561,
		24745	=>	55559,
		24746	=>	55557,
		24747	=>	55555,
		24748	=>	55552,
		24749	=>	55550,
		24750	=>	55548,
		24751	=>	55546,
		24752	=>	55543,
		24753	=>	55541,
		24754	=>	55539,
		24755	=>	55537,
		24756	=>	55534,
		24757	=>	55532,
		24758	=>	55530,
		24759	=>	55528,
		24760	=>	55525,
		24761	=>	55523,
		24762	=>	55521,
		24763	=>	55519,
		24764	=>	55516,
		24765	=>	55514,
		24766	=>	55512,
		24767	=>	55509,
		24768	=>	55507,
		24769	=>	55505,
		24770	=>	55503,
		24771	=>	55500,
		24772	=>	55498,
		24773	=>	55496,
		24774	=>	55494,
		24775	=>	55491,
		24776	=>	55489,
		24777	=>	55487,
		24778	=>	55485,
		24779	=>	55482,
		24780	=>	55480,
		24781	=>	55478,
		24782	=>	55476,
		24783	=>	55473,
		24784	=>	55471,
		24785	=>	55469,
		24786	=>	55466,
		24787	=>	55464,
		24788	=>	55462,
		24789	=>	55460,
		24790	=>	55457,
		24791	=>	55455,
		24792	=>	55453,
		24793	=>	55451,
		24794	=>	55448,
		24795	=>	55446,
		24796	=>	55444,
		24797	=>	55442,
		24798	=>	55439,
		24799	=>	55437,
		24800	=>	55435,
		24801	=>	55432,
		24802	=>	55430,
		24803	=>	55428,
		24804	=>	55426,
		24805	=>	55423,
		24806	=>	55421,
		24807	=>	55419,
		24808	=>	55417,
		24809	=>	55414,
		24810	=>	55412,
		24811	=>	55410,
		24812	=>	55407,
		24813	=>	55405,
		24814	=>	55403,
		24815	=>	55401,
		24816	=>	55398,
		24817	=>	55396,
		24818	=>	55394,
		24819	=>	55392,
		24820	=>	55389,
		24821	=>	55387,
		24822	=>	55385,
		24823	=>	55382,
		24824	=>	55380,
		24825	=>	55378,
		24826	=>	55376,
		24827	=>	55373,
		24828	=>	55371,
		24829	=>	55369,
		24830	=>	55367,
		24831	=>	55364,
		24832	=>	55362,
		24833	=>	55360,
		24834	=>	55357,
		24835	=>	55355,
		24836	=>	55353,
		24837	=>	55351,
		24838	=>	55348,
		24839	=>	55346,
		24840	=>	55344,
		24841	=>	55342,
		24842	=>	55339,
		24843	=>	55337,
		24844	=>	55335,
		24845	=>	55332,
		24846	=>	55330,
		24847	=>	55328,
		24848	=>	55326,
		24849	=>	55323,
		24850	=>	55321,
		24851	=>	55319,
		24852	=>	55316,
		24853	=>	55314,
		24854	=>	55312,
		24855	=>	55310,
		24856	=>	55307,
		24857	=>	55305,
		24858	=>	55303,
		24859	=>	55301,
		24860	=>	55298,
		24861	=>	55296,
		24862	=>	55294,
		24863	=>	55291,
		24864	=>	55289,
		24865	=>	55287,
		24866	=>	55285,
		24867	=>	55282,
		24868	=>	55280,
		24869	=>	55278,
		24870	=>	55275,
		24871	=>	55273,
		24872	=>	55271,
		24873	=>	55269,
		24874	=>	55266,
		24875	=>	55264,
		24876	=>	55262,
		24877	=>	55259,
		24878	=>	55257,
		24879	=>	55255,
		24880	=>	55253,
		24881	=>	55250,
		24882	=>	55248,
		24883	=>	55246,
		24884	=>	55243,
		24885	=>	55241,
		24886	=>	55239,
		24887	=>	55237,
		24888	=>	55234,
		24889	=>	55232,
		24890	=>	55230,
		24891	=>	55227,
		24892	=>	55225,
		24893	=>	55223,
		24894	=>	55221,
		24895	=>	55218,
		24896	=>	55216,
		24897	=>	55214,
		24898	=>	55211,
		24899	=>	55209,
		24900	=>	55207,
		24901	=>	55205,
		24902	=>	55202,
		24903	=>	55200,
		24904	=>	55198,
		24905	=>	55195,
		24906	=>	55193,
		24907	=>	55191,
		24908	=>	55189,
		24909	=>	55186,
		24910	=>	55184,
		24911	=>	55182,
		24912	=>	55179,
		24913	=>	55177,
		24914	=>	55175,
		24915	=>	55172,
		24916	=>	55170,
		24917	=>	55168,
		24918	=>	55166,
		24919	=>	55163,
		24920	=>	55161,
		24921	=>	55159,
		24922	=>	55156,
		24923	=>	55154,
		24924	=>	55152,
		24925	=>	55150,
		24926	=>	55147,
		24927	=>	55145,
		24928	=>	55143,
		24929	=>	55140,
		24930	=>	55138,
		24931	=>	55136,
		24932	=>	55133,
		24933	=>	55131,
		24934	=>	55129,
		24935	=>	55127,
		24936	=>	55124,
		24937	=>	55122,
		24938	=>	55120,
		24939	=>	55117,
		24940	=>	55115,
		24941	=>	55113,
		24942	=>	55110,
		24943	=>	55108,
		24944	=>	55106,
		24945	=>	55104,
		24946	=>	55101,
		24947	=>	55099,
		24948	=>	55097,
		24949	=>	55094,
		24950	=>	55092,
		24951	=>	55090,
		24952	=>	55087,
		24953	=>	55085,
		24954	=>	55083,
		24955	=>	55081,
		24956	=>	55078,
		24957	=>	55076,
		24958	=>	55074,
		24959	=>	55071,
		24960	=>	55069,
		24961	=>	55067,
		24962	=>	55064,
		24963	=>	55062,
		24964	=>	55060,
		24965	=>	55058,
		24966	=>	55055,
		24967	=>	55053,
		24968	=>	55051,
		24969	=>	55048,
		24970	=>	55046,
		24971	=>	55044,
		24972	=>	55041,
		24973	=>	55039,
		24974	=>	55037,
		24975	=>	55035,
		24976	=>	55032,
		24977	=>	55030,
		24978	=>	55028,
		24979	=>	55025,
		24980	=>	55023,
		24981	=>	55021,
		24982	=>	55018,
		24983	=>	55016,
		24984	=>	55014,
		24985	=>	55011,
		24986	=>	55009,
		24987	=>	55007,
		24988	=>	55005,
		24989	=>	55002,
		24990	=>	55000,
		24991	=>	54998,
		24992	=>	54995,
		24993	=>	54993,
		24994	=>	54991,
		24995	=>	54988,
		24996	=>	54986,
		24997	=>	54984,
		24998	=>	54981,
		24999	=>	54979,
		25000	=>	54977,
		25001	=>	54975,
		25002	=>	54972,
		25003	=>	54970,
		25004	=>	54968,
		25005	=>	54965,
		25006	=>	54963,
		25007	=>	54961,
		25008	=>	54958,
		25009	=>	54956,
		25010	=>	54954,
		25011	=>	54951,
		25012	=>	54949,
		25013	=>	54947,
		25014	=>	54945,
		25015	=>	54942,
		25016	=>	54940,
		25017	=>	54938,
		25018	=>	54935,
		25019	=>	54933,
		25020	=>	54931,
		25021	=>	54928,
		25022	=>	54926,
		25023	=>	54924,
		25024	=>	54921,
		25025	=>	54919,
		25026	=>	54917,
		25027	=>	54914,
		25028	=>	54912,
		25029	=>	54910,
		25030	=>	54907,
		25031	=>	54905,
		25032	=>	54903,
		25033	=>	54901,
		25034	=>	54898,
		25035	=>	54896,
		25036	=>	54894,
		25037	=>	54891,
		25038	=>	54889,
		25039	=>	54887,
		25040	=>	54884,
		25041	=>	54882,
		25042	=>	54880,
		25043	=>	54877,
		25044	=>	54875,
		25045	=>	54873,
		25046	=>	54870,
		25047	=>	54868,
		25048	=>	54866,
		25049	=>	54863,
		25050	=>	54861,
		25051	=>	54859,
		25052	=>	54856,
		25053	=>	54854,
		25054	=>	54852,
		25055	=>	54850,
		25056	=>	54847,
		25057	=>	54845,
		25058	=>	54843,
		25059	=>	54840,
		25060	=>	54838,
		25061	=>	54836,
		25062	=>	54833,
		25063	=>	54831,
		25064	=>	54829,
		25065	=>	54826,
		25066	=>	54824,
		25067	=>	54822,
		25068	=>	54819,
		25069	=>	54817,
		25070	=>	54815,
		25071	=>	54812,
		25072	=>	54810,
		25073	=>	54808,
		25074	=>	54805,
		25075	=>	54803,
		25076	=>	54801,
		25077	=>	54798,
		25078	=>	54796,
		25079	=>	54794,
		25080	=>	54791,
		25081	=>	54789,
		25082	=>	54787,
		25083	=>	54784,
		25084	=>	54782,
		25085	=>	54780,
		25086	=>	54777,
		25087	=>	54775,
		25088	=>	54773,
		25089	=>	54770,
		25090	=>	54768,
		25091	=>	54766,
		25092	=>	54763,
		25093	=>	54761,
		25094	=>	54759,
		25095	=>	54757,
		25096	=>	54754,
		25097	=>	54752,
		25098	=>	54750,
		25099	=>	54747,
		25100	=>	54745,
		25101	=>	54743,
		25102	=>	54740,
		25103	=>	54738,
		25104	=>	54736,
		25105	=>	54733,
		25106	=>	54731,
		25107	=>	54729,
		25108	=>	54726,
		25109	=>	54724,
		25110	=>	54722,
		25111	=>	54719,
		25112	=>	54717,
		25113	=>	54715,
		25114	=>	54712,
		25115	=>	54710,
		25116	=>	54708,
		25117	=>	54705,
		25118	=>	54703,
		25119	=>	54701,
		25120	=>	54698,
		25121	=>	54696,
		25122	=>	54694,
		25123	=>	54691,
		25124	=>	54689,
		25125	=>	54687,
		25126	=>	54684,
		25127	=>	54682,
		25128	=>	54680,
		25129	=>	54677,
		25130	=>	54675,
		25131	=>	54673,
		25132	=>	54670,
		25133	=>	54668,
		25134	=>	54666,
		25135	=>	54663,
		25136	=>	54661,
		25137	=>	54659,
		25138	=>	54656,
		25139	=>	54654,
		25140	=>	54651,
		25141	=>	54649,
		25142	=>	54647,
		25143	=>	54644,
		25144	=>	54642,
		25145	=>	54640,
		25146	=>	54637,
		25147	=>	54635,
		25148	=>	54633,
		25149	=>	54630,
		25150	=>	54628,
		25151	=>	54626,
		25152	=>	54623,
		25153	=>	54621,
		25154	=>	54619,
		25155	=>	54616,
		25156	=>	54614,
		25157	=>	54612,
		25158	=>	54609,
		25159	=>	54607,
		25160	=>	54605,
		25161	=>	54602,
		25162	=>	54600,
		25163	=>	54598,
		25164	=>	54595,
		25165	=>	54593,
		25166	=>	54591,
		25167	=>	54588,
		25168	=>	54586,
		25169	=>	54584,
		25170	=>	54581,
		25171	=>	54579,
		25172	=>	54577,
		25173	=>	54574,
		25174	=>	54572,
		25175	=>	54570,
		25176	=>	54567,
		25177	=>	54565,
		25178	=>	54562,
		25179	=>	54560,
		25180	=>	54558,
		25181	=>	54555,
		25182	=>	54553,
		25183	=>	54551,
		25184	=>	54548,
		25185	=>	54546,
		25186	=>	54544,
		25187	=>	54541,
		25188	=>	54539,
		25189	=>	54537,
		25190	=>	54534,
		25191	=>	54532,
		25192	=>	54530,
		25193	=>	54527,
		25194	=>	54525,
		25195	=>	54523,
		25196	=>	54520,
		25197	=>	54518,
		25198	=>	54516,
		25199	=>	54513,
		25200	=>	54511,
		25201	=>	54508,
		25202	=>	54506,
		25203	=>	54504,
		25204	=>	54501,
		25205	=>	54499,
		25206	=>	54497,
		25207	=>	54494,
		25208	=>	54492,
		25209	=>	54490,
		25210	=>	54487,
		25211	=>	54485,
		25212	=>	54483,
		25213	=>	54480,
		25214	=>	54478,
		25215	=>	54476,
		25216	=>	54473,
		25217	=>	54471,
		25218	=>	54469,
		25219	=>	54466,
		25220	=>	54464,
		25221	=>	54461,
		25222	=>	54459,
		25223	=>	54457,
		25224	=>	54454,
		25225	=>	54452,
		25226	=>	54450,
		25227	=>	54447,
		25228	=>	54445,
		25229	=>	54443,
		25230	=>	54440,
		25231	=>	54438,
		25232	=>	54436,
		25233	=>	54433,
		25234	=>	54431,
		25235	=>	54428,
		25236	=>	54426,
		25237	=>	54424,
		25238	=>	54421,
		25239	=>	54419,
		25240	=>	54417,
		25241	=>	54414,
		25242	=>	54412,
		25243	=>	54410,
		25244	=>	54407,
		25245	=>	54405,
		25246	=>	54403,
		25247	=>	54400,
		25248	=>	54398,
		25249	=>	54395,
		25250	=>	54393,
		25251	=>	54391,
		25252	=>	54388,
		25253	=>	54386,
		25254	=>	54384,
		25255	=>	54381,
		25256	=>	54379,
		25257	=>	54377,
		25258	=>	54374,
		25259	=>	54372,
		25260	=>	54369,
		25261	=>	54367,
		25262	=>	54365,
		25263	=>	54362,
		25264	=>	54360,
		25265	=>	54358,
		25266	=>	54355,
		25267	=>	54353,
		25268	=>	54351,
		25269	=>	54348,
		25270	=>	54346,
		25271	=>	54343,
		25272	=>	54341,
		25273	=>	54339,
		25274	=>	54336,
		25275	=>	54334,
		25276	=>	54332,
		25277	=>	54329,
		25278	=>	54327,
		25279	=>	54325,
		25280	=>	54322,
		25281	=>	54320,
		25282	=>	54317,
		25283	=>	54315,
		25284	=>	54313,
		25285	=>	54310,
		25286	=>	54308,
		25287	=>	54306,
		25288	=>	54303,
		25289	=>	54301,
		25290	=>	54299,
		25291	=>	54296,
		25292	=>	54294,
		25293	=>	54291,
		25294	=>	54289,
		25295	=>	54287,
		25296	=>	54284,
		25297	=>	54282,
		25298	=>	54280,
		25299	=>	54277,
		25300	=>	54275,
		25301	=>	54272,
		25302	=>	54270,
		25303	=>	54268,
		25304	=>	54265,
		25305	=>	54263,
		25306	=>	54261,
		25307	=>	54258,
		25308	=>	54256,
		25309	=>	54253,
		25310	=>	54251,
		25311	=>	54249,
		25312	=>	54246,
		25313	=>	54244,
		25314	=>	54242,
		25315	=>	54239,
		25316	=>	54237,
		25317	=>	54234,
		25318	=>	54232,
		25319	=>	54230,
		25320	=>	54227,
		25321	=>	54225,
		25322	=>	54223,
		25323	=>	54220,
		25324	=>	54218,
		25325	=>	54216,
		25326	=>	54213,
		25327	=>	54211,
		25328	=>	54208,
		25329	=>	54206,
		25330	=>	54204,
		25331	=>	54201,
		25332	=>	54199,
		25333	=>	54196,
		25334	=>	54194,
		25335	=>	54192,
		25336	=>	54189,
		25337	=>	54187,
		25338	=>	54185,
		25339	=>	54182,
		25340	=>	54180,
		25341	=>	54177,
		25342	=>	54175,
		25343	=>	54173,
		25344	=>	54170,
		25345	=>	54168,
		25346	=>	54166,
		25347	=>	54163,
		25348	=>	54161,
		25349	=>	54158,
		25350	=>	54156,
		25351	=>	54154,
		25352	=>	54151,
		25353	=>	54149,
		25354	=>	54147,
		25355	=>	54144,
		25356	=>	54142,
		25357	=>	54139,
		25358	=>	54137,
		25359	=>	54135,
		25360	=>	54132,
		25361	=>	54130,
		25362	=>	54127,
		25363	=>	54125,
		25364	=>	54123,
		25365	=>	54120,
		25366	=>	54118,
		25367	=>	54116,
		25368	=>	54113,
		25369	=>	54111,
		25370	=>	54108,
		25371	=>	54106,
		25372	=>	54104,
		25373	=>	54101,
		25374	=>	54099,
		25375	=>	54097,
		25376	=>	54094,
		25377	=>	54092,
		25378	=>	54089,
		25379	=>	54087,
		25380	=>	54085,
		25381	=>	54082,
		25382	=>	54080,
		25383	=>	54077,
		25384	=>	54075,
		25385	=>	54073,
		25386	=>	54070,
		25387	=>	54068,
		25388	=>	54065,
		25389	=>	54063,
		25390	=>	54061,
		25391	=>	54058,
		25392	=>	54056,
		25393	=>	54054,
		25394	=>	54051,
		25395	=>	54049,
		25396	=>	54046,
		25397	=>	54044,
		25398	=>	54042,
		25399	=>	54039,
		25400	=>	54037,
		25401	=>	54034,
		25402	=>	54032,
		25403	=>	54030,
		25404	=>	54027,
		25405	=>	54025,
		25406	=>	54022,
		25407	=>	54020,
		25408	=>	54018,
		25409	=>	54015,
		25410	=>	54013,
		25411	=>	54011,
		25412	=>	54008,
		25413	=>	54006,
		25414	=>	54003,
		25415	=>	54001,
		25416	=>	53999,
		25417	=>	53996,
		25418	=>	53994,
		25419	=>	53991,
		25420	=>	53989,
		25421	=>	53987,
		25422	=>	53984,
		25423	=>	53982,
		25424	=>	53979,
		25425	=>	53977,
		25426	=>	53975,
		25427	=>	53972,
		25428	=>	53970,
		25429	=>	53967,
		25430	=>	53965,
		25431	=>	53963,
		25432	=>	53960,
		25433	=>	53958,
		25434	=>	53955,
		25435	=>	53953,
		25436	=>	53951,
		25437	=>	53948,
		25438	=>	53946,
		25439	=>	53943,
		25440	=>	53941,
		25441	=>	53939,
		25442	=>	53936,
		25443	=>	53934,
		25444	=>	53931,
		25445	=>	53929,
		25446	=>	53927,
		25447	=>	53924,
		25448	=>	53922,
		25449	=>	53919,
		25450	=>	53917,
		25451	=>	53915,
		25452	=>	53912,
		25453	=>	53910,
		25454	=>	53907,
		25455	=>	53905,
		25456	=>	53903,
		25457	=>	53900,
		25458	=>	53898,
		25459	=>	53895,
		25460	=>	53893,
		25461	=>	53891,
		25462	=>	53888,
		25463	=>	53886,
		25464	=>	53883,
		25465	=>	53881,
		25466	=>	53879,
		25467	=>	53876,
		25468	=>	53874,
		25469	=>	53871,
		25470	=>	53869,
		25471	=>	53867,
		25472	=>	53864,
		25473	=>	53862,
		25474	=>	53859,
		25475	=>	53857,
		25476	=>	53855,
		25477	=>	53852,
		25478	=>	53850,
		25479	=>	53847,
		25480	=>	53845,
		25481	=>	53843,
		25482	=>	53840,
		25483	=>	53838,
		25484	=>	53835,
		25485	=>	53833,
		25486	=>	53831,
		25487	=>	53828,
		25488	=>	53826,
		25489	=>	53823,
		25490	=>	53821,
		25491	=>	53819,
		25492	=>	53816,
		25493	=>	53814,
		25494	=>	53811,
		25495	=>	53809,
		25496	=>	53807,
		25497	=>	53804,
		25498	=>	53802,
		25499	=>	53799,
		25500	=>	53797,
		25501	=>	53794,
		25502	=>	53792,
		25503	=>	53790,
		25504	=>	53787,
		25505	=>	53785,
		25506	=>	53782,
		25507	=>	53780,
		25508	=>	53778,
		25509	=>	53775,
		25510	=>	53773,
		25511	=>	53770,
		25512	=>	53768,
		25513	=>	53766,
		25514	=>	53763,
		25515	=>	53761,
		25516	=>	53758,
		25517	=>	53756,
		25518	=>	53753,
		25519	=>	53751,
		25520	=>	53749,
		25521	=>	53746,
		25522	=>	53744,
		25523	=>	53741,
		25524	=>	53739,
		25525	=>	53737,
		25526	=>	53734,
		25527	=>	53732,
		25528	=>	53729,
		25529	=>	53727,
		25530	=>	53725,
		25531	=>	53722,
		25532	=>	53720,
		25533	=>	53717,
		25534	=>	53715,
		25535	=>	53712,
		25536	=>	53710,
		25537	=>	53708,
		25538	=>	53705,
		25539	=>	53703,
		25540	=>	53700,
		25541	=>	53698,
		25542	=>	53696,
		25543	=>	53693,
		25544	=>	53691,
		25545	=>	53688,
		25546	=>	53686,
		25547	=>	53683,
		25548	=>	53681,
		25549	=>	53679,
		25550	=>	53676,
		25551	=>	53674,
		25552	=>	53671,
		25553	=>	53669,
		25554	=>	53666,
		25555	=>	53664,
		25556	=>	53662,
		25557	=>	53659,
		25558	=>	53657,
		25559	=>	53654,
		25560	=>	53652,
		25561	=>	53650,
		25562	=>	53647,
		25563	=>	53645,
		25564	=>	53642,
		25565	=>	53640,
		25566	=>	53637,
		25567	=>	53635,
		25568	=>	53633,
		25569	=>	53630,
		25570	=>	53628,
		25571	=>	53625,
		25572	=>	53623,
		25573	=>	53620,
		25574	=>	53618,
		25575	=>	53616,
		25576	=>	53613,
		25577	=>	53611,
		25578	=>	53608,
		25579	=>	53606,
		25580	=>	53604,
		25581	=>	53601,
		25582	=>	53599,
		25583	=>	53596,
		25584	=>	53594,
		25585	=>	53591,
		25586	=>	53589,
		25587	=>	53587,
		25588	=>	53584,
		25589	=>	53582,
		25590	=>	53579,
		25591	=>	53577,
		25592	=>	53574,
		25593	=>	53572,
		25594	=>	53570,
		25595	=>	53567,
		25596	=>	53565,
		25597	=>	53562,
		25598	=>	53560,
		25599	=>	53557,
		25600	=>	53555,
		25601	=>	53553,
		25602	=>	53550,
		25603	=>	53548,
		25604	=>	53545,
		25605	=>	53543,
		25606	=>	53540,
		25607	=>	53538,
		25608	=>	53536,
		25609	=>	53533,
		25610	=>	53531,
		25611	=>	53528,
		25612	=>	53526,
		25613	=>	53523,
		25614	=>	53521,
		25615	=>	53519,
		25616	=>	53516,
		25617	=>	53514,
		25618	=>	53511,
		25619	=>	53509,
		25620	=>	53506,
		25621	=>	53504,
		25622	=>	53502,
		25623	=>	53499,
		25624	=>	53497,
		25625	=>	53494,
		25626	=>	53492,
		25627	=>	53489,
		25628	=>	53487,
		25629	=>	53484,
		25630	=>	53482,
		25631	=>	53480,
		25632	=>	53477,
		25633	=>	53475,
		25634	=>	53472,
		25635	=>	53470,
		25636	=>	53467,
		25637	=>	53465,
		25638	=>	53463,
		25639	=>	53460,
		25640	=>	53458,
		25641	=>	53455,
		25642	=>	53453,
		25643	=>	53450,
		25644	=>	53448,
		25645	=>	53446,
		25646	=>	53443,
		25647	=>	53441,
		25648	=>	53438,
		25649	=>	53436,
		25650	=>	53433,
		25651	=>	53431,
		25652	=>	53428,
		25653	=>	53426,
		25654	=>	53424,
		25655	=>	53421,
		25656	=>	53419,
		25657	=>	53416,
		25658	=>	53414,
		25659	=>	53411,
		25660	=>	53409,
		25661	=>	53406,
		25662	=>	53404,
		25663	=>	53402,
		25664	=>	53399,
		25665	=>	53397,
		25666	=>	53394,
		25667	=>	53392,
		25668	=>	53389,
		25669	=>	53387,
		25670	=>	53385,
		25671	=>	53382,
		25672	=>	53380,
		25673	=>	53377,
		25674	=>	53375,
		25675	=>	53372,
		25676	=>	53370,
		25677	=>	53367,
		25678	=>	53365,
		25679	=>	53363,
		25680	=>	53360,
		25681	=>	53358,
		25682	=>	53355,
		25683	=>	53353,
		25684	=>	53350,
		25685	=>	53348,
		25686	=>	53345,
		25687	=>	53343,
		25688	=>	53341,
		25689	=>	53338,
		25690	=>	53336,
		25691	=>	53333,
		25692	=>	53331,
		25693	=>	53328,
		25694	=>	53326,
		25695	=>	53323,
		25696	=>	53321,
		25697	=>	53319,
		25698	=>	53316,
		25699	=>	53314,
		25700	=>	53311,
		25701	=>	53309,
		25702	=>	53306,
		25703	=>	53304,
		25704	=>	53301,
		25705	=>	53299,
		25706	=>	53296,
		25707	=>	53294,
		25708	=>	53292,
		25709	=>	53289,
		25710	=>	53287,
		25711	=>	53284,
		25712	=>	53282,
		25713	=>	53279,
		25714	=>	53277,
		25715	=>	53274,
		25716	=>	53272,
		25717	=>	53270,
		25718	=>	53267,
		25719	=>	53265,
		25720	=>	53262,
		25721	=>	53260,
		25722	=>	53257,
		25723	=>	53255,
		25724	=>	53252,
		25725	=>	53250,
		25726	=>	53247,
		25727	=>	53245,
		25728	=>	53243,
		25729	=>	53240,
		25730	=>	53238,
		25731	=>	53235,
		25732	=>	53233,
		25733	=>	53230,
		25734	=>	53228,
		25735	=>	53225,
		25736	=>	53223,
		25737	=>	53221,
		25738	=>	53218,
		25739	=>	53216,
		25740	=>	53213,
		25741	=>	53211,
		25742	=>	53208,
		25743	=>	53206,
		25744	=>	53203,
		25745	=>	53201,
		25746	=>	53198,
		25747	=>	53196,
		25748	=>	53193,
		25749	=>	53191,
		25750	=>	53189,
		25751	=>	53186,
		25752	=>	53184,
		25753	=>	53181,
		25754	=>	53179,
		25755	=>	53176,
		25756	=>	53174,
		25757	=>	53171,
		25758	=>	53169,
		25759	=>	53166,
		25760	=>	53164,
		25761	=>	53162,
		25762	=>	53159,
		25763	=>	53157,
		25764	=>	53154,
		25765	=>	53152,
		25766	=>	53149,
		25767	=>	53147,
		25768	=>	53144,
		25769	=>	53142,
		25770	=>	53139,
		25771	=>	53137,
		25772	=>	53134,
		25773	=>	53132,
		25774	=>	53130,
		25775	=>	53127,
		25776	=>	53125,
		25777	=>	53122,
		25778	=>	53120,
		25779	=>	53117,
		25780	=>	53115,
		25781	=>	53112,
		25782	=>	53110,
		25783	=>	53107,
		25784	=>	53105,
		25785	=>	53102,
		25786	=>	53100,
		25787	=>	53098,
		25788	=>	53095,
		25789	=>	53093,
		25790	=>	53090,
		25791	=>	53088,
		25792	=>	53085,
		25793	=>	53083,
		25794	=>	53080,
		25795	=>	53078,
		25796	=>	53075,
		25797	=>	53073,
		25798	=>	53070,
		25799	=>	53068,
		25800	=>	53066,
		25801	=>	53063,
		25802	=>	53061,
		25803	=>	53058,
		25804	=>	53056,
		25805	=>	53053,
		25806	=>	53051,
		25807	=>	53048,
		25808	=>	53046,
		25809	=>	53043,
		25810	=>	53041,
		25811	=>	53038,
		25812	=>	53036,
		25813	=>	53033,
		25814	=>	53031,
		25815	=>	53028,
		25816	=>	53026,
		25817	=>	53024,
		25818	=>	53021,
		25819	=>	53019,
		25820	=>	53016,
		25821	=>	53014,
		25822	=>	53011,
		25823	=>	53009,
		25824	=>	53006,
		25825	=>	53004,
		25826	=>	53001,
		25827	=>	52999,
		25828	=>	52996,
		25829	=>	52994,
		25830	=>	52991,
		25831	=>	52989,
		25832	=>	52986,
		25833	=>	52984,
		25834	=>	52982,
		25835	=>	52979,
		25836	=>	52977,
		25837	=>	52974,
		25838	=>	52972,
		25839	=>	52969,
		25840	=>	52967,
		25841	=>	52964,
		25842	=>	52962,
		25843	=>	52959,
		25844	=>	52957,
		25845	=>	52954,
		25846	=>	52952,
		25847	=>	52949,
		25848	=>	52947,
		25849	=>	52944,
		25850	=>	52942,
		25851	=>	52939,
		25852	=>	52937,
		25853	=>	52935,
		25854	=>	52932,
		25855	=>	52930,
		25856	=>	52927,
		25857	=>	52925,
		25858	=>	52922,
		25859	=>	52920,
		25860	=>	52917,
		25861	=>	52915,
		25862	=>	52912,
		25863	=>	52910,
		25864	=>	52907,
		25865	=>	52905,
		25866	=>	52902,
		25867	=>	52900,
		25868	=>	52897,
		25869	=>	52895,
		25870	=>	52892,
		25871	=>	52890,
		25872	=>	52887,
		25873	=>	52885,
		25874	=>	52882,
		25875	=>	52880,
		25876	=>	52878,
		25877	=>	52875,
		25878	=>	52873,
		25879	=>	52870,
		25880	=>	52868,
		25881	=>	52865,
		25882	=>	52863,
		25883	=>	52860,
		25884	=>	52858,
		25885	=>	52855,
		25886	=>	52853,
		25887	=>	52850,
		25888	=>	52848,
		25889	=>	52845,
		25890	=>	52843,
		25891	=>	52840,
		25892	=>	52838,
		25893	=>	52835,
		25894	=>	52833,
		25895	=>	52830,
		25896	=>	52828,
		25897	=>	52825,
		25898	=>	52823,
		25899	=>	52820,
		25900	=>	52818,
		25901	=>	52815,
		25902	=>	52813,
		25903	=>	52810,
		25904	=>	52808,
		25905	=>	52806,
		25906	=>	52803,
		25907	=>	52801,
		25908	=>	52798,
		25909	=>	52796,
		25910	=>	52793,
		25911	=>	52791,
		25912	=>	52788,
		25913	=>	52786,
		25914	=>	52783,
		25915	=>	52781,
		25916	=>	52778,
		25917	=>	52776,
		25918	=>	52773,
		25919	=>	52771,
		25920	=>	52768,
		25921	=>	52766,
		25922	=>	52763,
		25923	=>	52761,
		25924	=>	52758,
		25925	=>	52756,
		25926	=>	52753,
		25927	=>	52751,
		25928	=>	52748,
		25929	=>	52746,
		25930	=>	52743,
		25931	=>	52741,
		25932	=>	52738,
		25933	=>	52736,
		25934	=>	52733,
		25935	=>	52731,
		25936	=>	52728,
		25937	=>	52726,
		25938	=>	52723,
		25939	=>	52721,
		25940	=>	52718,
		25941	=>	52716,
		25942	=>	52713,
		25943	=>	52711,
		25944	=>	52708,
		25945	=>	52706,
		25946	=>	52703,
		25947	=>	52701,
		25948	=>	52698,
		25949	=>	52696,
		25950	=>	52693,
		25951	=>	52691,
		25952	=>	52688,
		25953	=>	52686,
		25954	=>	52684,
		25955	=>	52681,
		25956	=>	52679,
		25957	=>	52676,
		25958	=>	52674,
		25959	=>	52671,
		25960	=>	52669,
		25961	=>	52666,
		25962	=>	52664,
		25963	=>	52661,
		25964	=>	52659,
		25965	=>	52656,
		25966	=>	52654,
		25967	=>	52651,
		25968	=>	52649,
		25969	=>	52646,
		25970	=>	52644,
		25971	=>	52641,
		25972	=>	52639,
		25973	=>	52636,
		25974	=>	52634,
		25975	=>	52631,
		25976	=>	52629,
		25977	=>	52626,
		25978	=>	52624,
		25979	=>	52621,
		25980	=>	52619,
		25981	=>	52616,
		25982	=>	52614,
		25983	=>	52611,
		25984	=>	52609,
		25985	=>	52606,
		25986	=>	52604,
		25987	=>	52601,
		25988	=>	52599,
		25989	=>	52596,
		25990	=>	52594,
		25991	=>	52591,
		25992	=>	52589,
		25993	=>	52586,
		25994	=>	52584,
		25995	=>	52581,
		25996	=>	52579,
		25997	=>	52576,
		25998	=>	52574,
		25999	=>	52571,
		26000	=>	52569,
		26001	=>	52566,
		26002	=>	52564,
		26003	=>	52561,
		26004	=>	52559,
		26005	=>	52556,
		26006	=>	52554,
		26007	=>	52551,
		26008	=>	52549,
		26009	=>	52546,
		26010	=>	52544,
		26011	=>	52541,
		26012	=>	52539,
		26013	=>	52536,
		26014	=>	52533,
		26015	=>	52531,
		26016	=>	52528,
		26017	=>	52526,
		26018	=>	52523,
		26019	=>	52521,
		26020	=>	52518,
		26021	=>	52516,
		26022	=>	52513,
		26023	=>	52511,
		26024	=>	52508,
		26025	=>	52506,
		26026	=>	52503,
		26027	=>	52501,
		26028	=>	52498,
		26029	=>	52496,
		26030	=>	52493,
		26031	=>	52491,
		26032	=>	52488,
		26033	=>	52486,
		26034	=>	52483,
		26035	=>	52481,
		26036	=>	52478,
		26037	=>	52476,
		26038	=>	52473,
		26039	=>	52471,
		26040	=>	52468,
		26041	=>	52466,
		26042	=>	52463,
		26043	=>	52461,
		26044	=>	52458,
		26045	=>	52456,
		26046	=>	52453,
		26047	=>	52451,
		26048	=>	52448,
		26049	=>	52446,
		26050	=>	52443,
		26051	=>	52441,
		26052	=>	52438,
		26053	=>	52436,
		26054	=>	52433,
		26055	=>	52431,
		26056	=>	52428,
		26057	=>	52426,
		26058	=>	52423,
		26059	=>	52421,
		26060	=>	52418,
		26061	=>	52416,
		26062	=>	52413,
		26063	=>	52411,
		26064	=>	52408,
		26065	=>	52405,
		26066	=>	52403,
		26067	=>	52400,
		26068	=>	52398,
		26069	=>	52395,
		26070	=>	52393,
		26071	=>	52390,
		26072	=>	52388,
		26073	=>	52385,
		26074	=>	52383,
		26075	=>	52380,
		26076	=>	52378,
		26077	=>	52375,
		26078	=>	52373,
		26079	=>	52370,
		26080	=>	52368,
		26081	=>	52365,
		26082	=>	52363,
		26083	=>	52360,
		26084	=>	52358,
		26085	=>	52355,
		26086	=>	52353,
		26087	=>	52350,
		26088	=>	52348,
		26089	=>	52345,
		26090	=>	52343,
		26091	=>	52340,
		26092	=>	52338,
		26093	=>	52335,
		26094	=>	52332,
		26095	=>	52330,
		26096	=>	52327,
		26097	=>	52325,
		26098	=>	52322,
		26099	=>	52320,
		26100	=>	52317,
		26101	=>	52315,
		26102	=>	52312,
		26103	=>	52310,
		26104	=>	52307,
		26105	=>	52305,
		26106	=>	52302,
		26107	=>	52300,
		26108	=>	52297,
		26109	=>	52295,
		26110	=>	52292,
		26111	=>	52290,
		26112	=>	52287,
		26113	=>	52285,
		26114	=>	52282,
		26115	=>	52280,
		26116	=>	52277,
		26117	=>	52274,
		26118	=>	52272,
		26119	=>	52269,
		26120	=>	52267,
		26121	=>	52264,
		26122	=>	52262,
		26123	=>	52259,
		26124	=>	52257,
		26125	=>	52254,
		26126	=>	52252,
		26127	=>	52249,
		26128	=>	52247,
		26129	=>	52244,
		26130	=>	52242,
		26131	=>	52239,
		26132	=>	52237,
		26133	=>	52234,
		26134	=>	52232,
		26135	=>	52229,
		26136	=>	52226,
		26137	=>	52224,
		26138	=>	52221,
		26139	=>	52219,
		26140	=>	52216,
		26141	=>	52214,
		26142	=>	52211,
		26143	=>	52209,
		26144	=>	52206,
		26145	=>	52204,
		26146	=>	52201,
		26147	=>	52199,
		26148	=>	52196,
		26149	=>	52194,
		26150	=>	52191,
		26151	=>	52189,
		26152	=>	52186,
		26153	=>	52183,
		26154	=>	52181,
		26155	=>	52178,
		26156	=>	52176,
		26157	=>	52173,
		26158	=>	52171,
		26159	=>	52168,
		26160	=>	52166,
		26161	=>	52163,
		26162	=>	52161,
		26163	=>	52158,
		26164	=>	52156,
		26165	=>	52153,
		26166	=>	52151,
		26167	=>	52148,
		26168	=>	52145,
		26169	=>	52143,
		26170	=>	52140,
		26171	=>	52138,
		26172	=>	52135,
		26173	=>	52133,
		26174	=>	52130,
		26175	=>	52128,
		26176	=>	52125,
		26177	=>	52123,
		26178	=>	52120,
		26179	=>	52118,
		26180	=>	52115,
		26181	=>	52113,
		26182	=>	52110,
		26183	=>	52107,
		26184	=>	52105,
		26185	=>	52102,
		26186	=>	52100,
		26187	=>	52097,
		26188	=>	52095,
		26189	=>	52092,
		26190	=>	52090,
		26191	=>	52087,
		26192	=>	52085,
		26193	=>	52082,
		26194	=>	52080,
		26195	=>	52077,
		26196	=>	52074,
		26197	=>	52072,
		26198	=>	52069,
		26199	=>	52067,
		26200	=>	52064,
		26201	=>	52062,
		26202	=>	52059,
		26203	=>	52057,
		26204	=>	52054,
		26205	=>	52052,
		26206	=>	52049,
		26207	=>	52047,
		26208	=>	52044,
		26209	=>	52041,
		26210	=>	52039,
		26211	=>	52036,
		26212	=>	52034,
		26213	=>	52031,
		26214	=>	52029,
		26215	=>	52026,
		26216	=>	52024,
		26217	=>	52021,
		26218	=>	52019,
		26219	=>	52016,
		26220	=>	52014,
		26221	=>	52011,
		26222	=>	52008,
		26223	=>	52006,
		26224	=>	52003,
		26225	=>	52001,
		26226	=>	51998,
		26227	=>	51996,
		26228	=>	51993,
		26229	=>	51991,
		26230	=>	51988,
		26231	=>	51986,
		26232	=>	51983,
		26233	=>	51980,
		26234	=>	51978,
		26235	=>	51975,
		26236	=>	51973,
		26237	=>	51970,
		26238	=>	51968,
		26239	=>	51965,
		26240	=>	51963,
		26241	=>	51960,
		26242	=>	51958,
		26243	=>	51955,
		26244	=>	51952,
		26245	=>	51950,
		26246	=>	51947,
		26247	=>	51945,
		26248	=>	51942,
		26249	=>	51940,
		26250	=>	51937,
		26251	=>	51935,
		26252	=>	51932,
		26253	=>	51930,
		26254	=>	51927,
		26255	=>	51924,
		26256	=>	51922,
		26257	=>	51919,
		26258	=>	51917,
		26259	=>	51914,
		26260	=>	51912,
		26261	=>	51909,
		26262	=>	51907,
		26263	=>	51904,
		26264	=>	51901,
		26265	=>	51899,
		26266	=>	51896,
		26267	=>	51894,
		26268	=>	51891,
		26269	=>	51889,
		26270	=>	51886,
		26271	=>	51884,
		26272	=>	51881,
		26273	=>	51879,
		26274	=>	51876,
		26275	=>	51873,
		26276	=>	51871,
		26277	=>	51868,
		26278	=>	51866,
		26279	=>	51863,
		26280	=>	51861,
		26281	=>	51858,
		26282	=>	51856,
		26283	=>	51853,
		26284	=>	51850,
		26285	=>	51848,
		26286	=>	51845,
		26287	=>	51843,
		26288	=>	51840,
		26289	=>	51838,
		26290	=>	51835,
		26291	=>	51833,
		26292	=>	51830,
		26293	=>	51827,
		26294	=>	51825,
		26295	=>	51822,
		26296	=>	51820,
		26297	=>	51817,
		26298	=>	51815,
		26299	=>	51812,
		26300	=>	51810,
		26301	=>	51807,
		26302	=>	51804,
		26303	=>	51802,
		26304	=>	51799,
		26305	=>	51797,
		26306	=>	51794,
		26307	=>	51792,
		26308	=>	51789,
		26309	=>	51787,
		26310	=>	51784,
		26311	=>	51781,
		26312	=>	51779,
		26313	=>	51776,
		26314	=>	51774,
		26315	=>	51771,
		26316	=>	51769,
		26317	=>	51766,
		26318	=>	51764,
		26319	=>	51761,
		26320	=>	51758,
		26321	=>	51756,
		26322	=>	51753,
		26323	=>	51751,
		26324	=>	51748,
		26325	=>	51746,
		26326	=>	51743,
		26327	=>	51740,
		26328	=>	51738,
		26329	=>	51735,
		26330	=>	51733,
		26331	=>	51730,
		26332	=>	51728,
		26333	=>	51725,
		26334	=>	51723,
		26335	=>	51720,
		26336	=>	51717,
		26337	=>	51715,
		26338	=>	51712,
		26339	=>	51710,
		26340	=>	51707,
		26341	=>	51705,
		26342	=>	51702,
		26343	=>	51699,
		26344	=>	51697,
		26345	=>	51694,
		26346	=>	51692,
		26347	=>	51689,
		26348	=>	51687,
		26349	=>	51684,
		26350	=>	51681,
		26351	=>	51679,
		26352	=>	51676,
		26353	=>	51674,
		26354	=>	51671,
		26355	=>	51669,
		26356	=>	51666,
		26357	=>	51664,
		26358	=>	51661,
		26359	=>	51658,
		26360	=>	51656,
		26361	=>	51653,
		26362	=>	51651,
		26363	=>	51648,
		26364	=>	51646,
		26365	=>	51643,
		26366	=>	51640,
		26367	=>	51638,
		26368	=>	51635,
		26369	=>	51633,
		26370	=>	51630,
		26371	=>	51628,
		26372	=>	51625,
		26373	=>	51622,
		26374	=>	51620,
		26375	=>	51617,
		26376	=>	51615,
		26377	=>	51612,
		26378	=>	51610,
		26379	=>	51607,
		26380	=>	51604,
		26381	=>	51602,
		26382	=>	51599,
		26383	=>	51597,
		26384	=>	51594,
		26385	=>	51592,
		26386	=>	51589,
		26387	=>	51586,
		26388	=>	51584,
		26389	=>	51581,
		26390	=>	51579,
		26391	=>	51576,
		26392	=>	51574,
		26393	=>	51571,
		26394	=>	51568,
		26395	=>	51566,
		26396	=>	51563,
		26397	=>	51561,
		26398	=>	51558,
		26399	=>	51556,
		26400	=>	51553,
		26401	=>	51550,
		26402	=>	51548,
		26403	=>	51545,
		26404	=>	51543,
		26405	=>	51540,
		26406	=>	51538,
		26407	=>	51535,
		26408	=>	51532,
		26409	=>	51530,
		26410	=>	51527,
		26411	=>	51525,
		26412	=>	51522,
		26413	=>	51520,
		26414	=>	51517,
		26415	=>	51514,
		26416	=>	51512,
		26417	=>	51509,
		26418	=>	51507,
		26419	=>	51504,
		26420	=>	51502,
		26421	=>	51499,
		26422	=>	51496,
		26423	=>	51494,
		26424	=>	51491,
		26425	=>	51489,
		26426	=>	51486,
		26427	=>	51483,
		26428	=>	51481,
		26429	=>	51478,
		26430	=>	51476,
		26431	=>	51473,
		26432	=>	51471,
		26433	=>	51468,
		26434	=>	51465,
		26435	=>	51463,
		26436	=>	51460,
		26437	=>	51458,
		26438	=>	51455,
		26439	=>	51452,
		26440	=>	51450,
		26441	=>	51447,
		26442	=>	51445,
		26443	=>	51442,
		26444	=>	51440,
		26445	=>	51437,
		26446	=>	51434,
		26447	=>	51432,
		26448	=>	51429,
		26449	=>	51427,
		26450	=>	51424,
		26451	=>	51422,
		26452	=>	51419,
		26453	=>	51416,
		26454	=>	51414,
		26455	=>	51411,
		26456	=>	51409,
		26457	=>	51406,
		26458	=>	51403,
		26459	=>	51401,
		26460	=>	51398,
		26461	=>	51396,
		26462	=>	51393,
		26463	=>	51391,
		26464	=>	51388,
		26465	=>	51385,
		26466	=>	51383,
		26467	=>	51380,
		26468	=>	51378,
		26469	=>	51375,
		26470	=>	51372,
		26471	=>	51370,
		26472	=>	51367,
		26473	=>	51365,
		26474	=>	51362,
		26475	=>	51359,
		26476	=>	51357,
		26477	=>	51354,
		26478	=>	51352,
		26479	=>	51349,
		26480	=>	51347,
		26481	=>	51344,
		26482	=>	51341,
		26483	=>	51339,
		26484	=>	51336,
		26485	=>	51334,
		26486	=>	51331,
		26487	=>	51328,
		26488	=>	51326,
		26489	=>	51323,
		26490	=>	51321,
		26491	=>	51318,
		26492	=>	51315,
		26493	=>	51313,
		26494	=>	51310,
		26495	=>	51308,
		26496	=>	51305,
		26497	=>	51303,
		26498	=>	51300,
		26499	=>	51297,
		26500	=>	51295,
		26501	=>	51292,
		26502	=>	51290,
		26503	=>	51287,
		26504	=>	51284,
		26505	=>	51282,
		26506	=>	51279,
		26507	=>	51277,
		26508	=>	51274,
		26509	=>	51271,
		26510	=>	51269,
		26511	=>	51266,
		26512	=>	51264,
		26513	=>	51261,
		26514	=>	51258,
		26515	=>	51256,
		26516	=>	51253,
		26517	=>	51251,
		26518	=>	51248,
		26519	=>	51245,
		26520	=>	51243,
		26521	=>	51240,
		26522	=>	51238,
		26523	=>	51235,
		26524	=>	51233,
		26525	=>	51230,
		26526	=>	51227,
		26527	=>	51225,
		26528	=>	51222,
		26529	=>	51220,
		26530	=>	51217,
		26531	=>	51214,
		26532	=>	51212,
		26533	=>	51209,
		26534	=>	51207,
		26535	=>	51204,
		26536	=>	51201,
		26537	=>	51199,
		26538	=>	51196,
		26539	=>	51194,
		26540	=>	51191,
		26541	=>	51188,
		26542	=>	51186,
		26543	=>	51183,
		26544	=>	51181,
		26545	=>	51178,
		26546	=>	51175,
		26547	=>	51173,
		26548	=>	51170,
		26549	=>	51168,
		26550	=>	51165,
		26551	=>	51162,
		26552	=>	51160,
		26553	=>	51157,
		26554	=>	51155,
		26555	=>	51152,
		26556	=>	51149,
		26557	=>	51147,
		26558	=>	51144,
		26559	=>	51142,
		26560	=>	51139,
		26561	=>	51136,
		26562	=>	51134,
		26563	=>	51131,
		26564	=>	51129,
		26565	=>	51126,
		26566	=>	51123,
		26567	=>	51121,
		26568	=>	51118,
		26569	=>	51116,
		26570	=>	51113,
		26571	=>	51110,
		26572	=>	51108,
		26573	=>	51105,
		26574	=>	51103,
		26575	=>	51100,
		26576	=>	51097,
		26577	=>	51095,
		26578	=>	51092,
		26579	=>	51090,
		26580	=>	51087,
		26581	=>	51084,
		26582	=>	51082,
		26583	=>	51079,
		26584	=>	51076,
		26585	=>	51074,
		26586	=>	51071,
		26587	=>	51069,
		26588	=>	51066,
		26589	=>	51063,
		26590	=>	51061,
		26591	=>	51058,
		26592	=>	51056,
		26593	=>	51053,
		26594	=>	51050,
		26595	=>	51048,
		26596	=>	51045,
		26597	=>	51043,
		26598	=>	51040,
		26599	=>	51037,
		26600	=>	51035,
		26601	=>	51032,
		26602	=>	51030,
		26603	=>	51027,
		26604	=>	51024,
		26605	=>	51022,
		26606	=>	51019,
		26607	=>	51017,
		26608	=>	51014,
		26609	=>	51011,
		26610	=>	51009,
		26611	=>	51006,
		26612	=>	51003,
		26613	=>	51001,
		26614	=>	50998,
		26615	=>	50996,
		26616	=>	50993,
		26617	=>	50990,
		26618	=>	50988,
		26619	=>	50985,
		26620	=>	50983,
		26621	=>	50980,
		26622	=>	50977,
		26623	=>	50975,
		26624	=>	50972,
		26625	=>	50970,
		26626	=>	50967,
		26627	=>	50964,
		26628	=>	50962,
		26629	=>	50959,
		26630	=>	50956,
		26631	=>	50954,
		26632	=>	50951,
		26633	=>	50949,
		26634	=>	50946,
		26635	=>	50943,
		26636	=>	50941,
		26637	=>	50938,
		26638	=>	50936,
		26639	=>	50933,
		26640	=>	50930,
		26641	=>	50928,
		26642	=>	50925,
		26643	=>	50922,
		26644	=>	50920,
		26645	=>	50917,
		26646	=>	50915,
		26647	=>	50912,
		26648	=>	50909,
		26649	=>	50907,
		26650	=>	50904,
		26651	=>	50902,
		26652	=>	50899,
		26653	=>	50896,
		26654	=>	50894,
		26655	=>	50891,
		26656	=>	50888,
		26657	=>	50886,
		26658	=>	50883,
		26659	=>	50881,
		26660	=>	50878,
		26661	=>	50875,
		26662	=>	50873,
		26663	=>	50870,
		26664	=>	50868,
		26665	=>	50865,
		26666	=>	50862,
		26667	=>	50860,
		26668	=>	50857,
		26669	=>	50854,
		26670	=>	50852,
		26671	=>	50849,
		26672	=>	50847,
		26673	=>	50844,
		26674	=>	50841,
		26675	=>	50839,
		26676	=>	50836,
		26677	=>	50833,
		26678	=>	50831,
		26679	=>	50828,
		26680	=>	50826,
		26681	=>	50823,
		26682	=>	50820,
		26683	=>	50818,
		26684	=>	50815,
		26685	=>	50812,
		26686	=>	50810,
		26687	=>	50807,
		26688	=>	50805,
		26689	=>	50802,
		26690	=>	50799,
		26691	=>	50797,
		26692	=>	50794,
		26693	=>	50792,
		26694	=>	50789,
		26695	=>	50786,
		26696	=>	50784,
		26697	=>	50781,
		26698	=>	50778,
		26699	=>	50776,
		26700	=>	50773,
		26701	=>	50771,
		26702	=>	50768,
		26703	=>	50765,
		26704	=>	50763,
		26705	=>	50760,
		26706	=>	50757,
		26707	=>	50755,
		26708	=>	50752,
		26709	=>	50750,
		26710	=>	50747,
		26711	=>	50744,
		26712	=>	50742,
		26713	=>	50739,
		26714	=>	50736,
		26715	=>	50734,
		26716	=>	50731,
		26717	=>	50729,
		26718	=>	50726,
		26719	=>	50723,
		26720	=>	50721,
		26721	=>	50718,
		26722	=>	50715,
		26723	=>	50713,
		26724	=>	50710,
		26725	=>	50707,
		26726	=>	50705,
		26727	=>	50702,
		26728	=>	50700,
		26729	=>	50697,
		26730	=>	50694,
		26731	=>	50692,
		26732	=>	50689,
		26733	=>	50686,
		26734	=>	50684,
		26735	=>	50681,
		26736	=>	50679,
		26737	=>	50676,
		26738	=>	50673,
		26739	=>	50671,
		26740	=>	50668,
		26741	=>	50665,
		26742	=>	50663,
		26743	=>	50660,
		26744	=>	50657,
		26745	=>	50655,
		26746	=>	50652,
		26747	=>	50650,
		26748	=>	50647,
		26749	=>	50644,
		26750	=>	50642,
		26751	=>	50639,
		26752	=>	50636,
		26753	=>	50634,
		26754	=>	50631,
		26755	=>	50629,
		26756	=>	50626,
		26757	=>	50623,
		26758	=>	50621,
		26759	=>	50618,
		26760	=>	50615,
		26761	=>	50613,
		26762	=>	50610,
		26763	=>	50607,
		26764	=>	50605,
		26765	=>	50602,
		26766	=>	50600,
		26767	=>	50597,
		26768	=>	50594,
		26769	=>	50592,
		26770	=>	50589,
		26771	=>	50586,
		26772	=>	50584,
		26773	=>	50581,
		26774	=>	50578,
		26775	=>	50576,
		26776	=>	50573,
		26777	=>	50571,
		26778	=>	50568,
		26779	=>	50565,
		26780	=>	50563,
		26781	=>	50560,
		26782	=>	50557,
		26783	=>	50555,
		26784	=>	50552,
		26785	=>	50549,
		26786	=>	50547,
		26787	=>	50544,
		26788	=>	50542,
		26789	=>	50539,
		26790	=>	50536,
		26791	=>	50534,
		26792	=>	50531,
		26793	=>	50528,
		26794	=>	50526,
		26795	=>	50523,
		26796	=>	50520,
		26797	=>	50518,
		26798	=>	50515,
		26799	=>	50512,
		26800	=>	50510,
		26801	=>	50507,
		26802	=>	50505,
		26803	=>	50502,
		26804	=>	50499,
		26805	=>	50497,
		26806	=>	50494,
		26807	=>	50491,
		26808	=>	50489,
		26809	=>	50486,
		26810	=>	50483,
		26811	=>	50481,
		26812	=>	50478,
		26813	=>	50475,
		26814	=>	50473,
		26815	=>	50470,
		26816	=>	50468,
		26817	=>	50465,
		26818	=>	50462,
		26819	=>	50460,
		26820	=>	50457,
		26821	=>	50454,
		26822	=>	50452,
		26823	=>	50449,
		26824	=>	50446,
		26825	=>	50444,
		26826	=>	50441,
		26827	=>	50438,
		26828	=>	50436,
		26829	=>	50433,
		26830	=>	50431,
		26831	=>	50428,
		26832	=>	50425,
		26833	=>	50423,
		26834	=>	50420,
		26835	=>	50417,
		26836	=>	50415,
		26837	=>	50412,
		26838	=>	50409,
		26839	=>	50407,
		26840	=>	50404,
		26841	=>	50401,
		26842	=>	50399,
		26843	=>	50396,
		26844	=>	50393,
		26845	=>	50391,
		26846	=>	50388,
		26847	=>	50386,
		26848	=>	50383,
		26849	=>	50380,
		26850	=>	50378,
		26851	=>	50375,
		26852	=>	50372,
		26853	=>	50370,
		26854	=>	50367,
		26855	=>	50364,
		26856	=>	50362,
		26857	=>	50359,
		26858	=>	50356,
		26859	=>	50354,
		26860	=>	50351,
		26861	=>	50348,
		26862	=>	50346,
		26863	=>	50343,
		26864	=>	50340,
		26865	=>	50338,
		26866	=>	50335,
		26867	=>	50333,
		26868	=>	50330,
		26869	=>	50327,
		26870	=>	50325,
		26871	=>	50322,
		26872	=>	50319,
		26873	=>	50317,
		26874	=>	50314,
		26875	=>	50311,
		26876	=>	50309,
		26877	=>	50306,
		26878	=>	50303,
		26879	=>	50301,
		26880	=>	50298,
		26881	=>	50295,
		26882	=>	50293,
		26883	=>	50290,
		26884	=>	50287,
		26885	=>	50285,
		26886	=>	50282,
		26887	=>	50279,
		26888	=>	50277,
		26889	=>	50274,
		26890	=>	50271,
		26891	=>	50269,
		26892	=>	50266,
		26893	=>	50264,
		26894	=>	50261,
		26895	=>	50258,
		26896	=>	50256,
		26897	=>	50253,
		26898	=>	50250,
		26899	=>	50248,
		26900	=>	50245,
		26901	=>	50242,
		26902	=>	50240,
		26903	=>	50237,
		26904	=>	50234,
		26905	=>	50232,
		26906	=>	50229,
		26907	=>	50226,
		26908	=>	50224,
		26909	=>	50221,
		26910	=>	50218,
		26911	=>	50216,
		26912	=>	50213,
		26913	=>	50210,
		26914	=>	50208,
		26915	=>	50205,
		26916	=>	50202,
		26917	=>	50200,
		26918	=>	50197,
		26919	=>	50194,
		26920	=>	50192,
		26921	=>	50189,
		26922	=>	50186,
		26923	=>	50184,
		26924	=>	50181,
		26925	=>	50178,
		26926	=>	50176,
		26927	=>	50173,
		26928	=>	50170,
		26929	=>	50168,
		26930	=>	50165,
		26931	=>	50162,
		26932	=>	50160,
		26933	=>	50157,
		26934	=>	50154,
		26935	=>	50152,
		26936	=>	50149,
		26937	=>	50146,
		26938	=>	50144,
		26939	=>	50141,
		26940	=>	50138,
		26941	=>	50136,
		26942	=>	50133,
		26943	=>	50131,
		26944	=>	50128,
		26945	=>	50125,
		26946	=>	50123,
		26947	=>	50120,
		26948	=>	50117,
		26949	=>	50115,
		26950	=>	50112,
		26951	=>	50109,
		26952	=>	50107,
		26953	=>	50104,
		26954	=>	50101,
		26955	=>	50099,
		26956	=>	50096,
		26957	=>	50093,
		26958	=>	50091,
		26959	=>	50088,
		26960	=>	50085,
		26961	=>	50083,
		26962	=>	50080,
		26963	=>	50077,
		26964	=>	50075,
		26965	=>	50072,
		26966	=>	50069,
		26967	=>	50067,
		26968	=>	50064,
		26969	=>	50061,
		26970	=>	50059,
		26971	=>	50056,
		26972	=>	50053,
		26973	=>	50051,
		26974	=>	50048,
		26975	=>	50045,
		26976	=>	50042,
		26977	=>	50040,
		26978	=>	50037,
		26979	=>	50034,
		26980	=>	50032,
		26981	=>	50029,
		26982	=>	50026,
		26983	=>	50024,
		26984	=>	50021,
		26985	=>	50018,
		26986	=>	50016,
		26987	=>	50013,
		26988	=>	50010,
		26989	=>	50008,
		26990	=>	50005,
		26991	=>	50002,
		26992	=>	50000,
		26993	=>	49997,
		26994	=>	49994,
		26995	=>	49992,
		26996	=>	49989,
		26997	=>	49986,
		26998	=>	49984,
		26999	=>	49981,
		27000	=>	49978,
		27001	=>	49976,
		27002	=>	49973,
		27003	=>	49970,
		27004	=>	49968,
		27005	=>	49965,
		27006	=>	49962,
		27007	=>	49960,
		27008	=>	49957,
		27009	=>	49954,
		27010	=>	49952,
		27011	=>	49949,
		27012	=>	49946,
		27013	=>	49944,
		27014	=>	49941,
		27015	=>	49938,
		27016	=>	49936,
		27017	=>	49933,
		27018	=>	49930,
		27019	=>	49928,
		27020	=>	49925,
		27021	=>	49922,
		27022	=>	49920,
		27023	=>	49917,
		27024	=>	49914,
		27025	=>	49912,
		27026	=>	49909,
		27027	=>	49906,
		27028	=>	49903,
		27029	=>	49901,
		27030	=>	49898,
		27031	=>	49895,
		27032	=>	49893,
		27033	=>	49890,
		27034	=>	49887,
		27035	=>	49885,
		27036	=>	49882,
		27037	=>	49879,
		27038	=>	49877,
		27039	=>	49874,
		27040	=>	49871,
		27041	=>	49869,
		27042	=>	49866,
		27043	=>	49863,
		27044	=>	49861,
		27045	=>	49858,
		27046	=>	49855,
		27047	=>	49853,
		27048	=>	49850,
		27049	=>	49847,
		27050	=>	49845,
		27051	=>	49842,
		27052	=>	49839,
		27053	=>	49836,
		27054	=>	49834,
		27055	=>	49831,
		27056	=>	49828,
		27057	=>	49826,
		27058	=>	49823,
		27059	=>	49820,
		27060	=>	49818,
		27061	=>	49815,
		27062	=>	49812,
		27063	=>	49810,
		27064	=>	49807,
		27065	=>	49804,
		27066	=>	49802,
		27067	=>	49799,
		27068	=>	49796,
		27069	=>	49794,
		27070	=>	49791,
		27071	=>	49788,
		27072	=>	49785,
		27073	=>	49783,
		27074	=>	49780,
		27075	=>	49777,
		27076	=>	49775,
		27077	=>	49772,
		27078	=>	49769,
		27079	=>	49767,
		27080	=>	49764,
		27081	=>	49761,
		27082	=>	49759,
		27083	=>	49756,
		27084	=>	49753,
		27085	=>	49751,
		27086	=>	49748,
		27087	=>	49745,
		27088	=>	49743,
		27089	=>	49740,
		27090	=>	49737,
		27091	=>	49734,
		27092	=>	49732,
		27093	=>	49729,
		27094	=>	49726,
		27095	=>	49724,
		27096	=>	49721,
		27097	=>	49718,
		27098	=>	49716,
		27099	=>	49713,
		27100	=>	49710,
		27101	=>	49708,
		27102	=>	49705,
		27103	=>	49702,
		27104	=>	49700,
		27105	=>	49697,
		27106	=>	49694,
		27107	=>	49691,
		27108	=>	49689,
		27109	=>	49686,
		27110	=>	49683,
		27111	=>	49681,
		27112	=>	49678,
		27113	=>	49675,
		27114	=>	49673,
		27115	=>	49670,
		27116	=>	49667,
		27117	=>	49665,
		27118	=>	49662,
		27119	=>	49659,
		27120	=>	49656,
		27121	=>	49654,
		27122	=>	49651,
		27123	=>	49648,
		27124	=>	49646,
		27125	=>	49643,
		27126	=>	49640,
		27127	=>	49638,
		27128	=>	49635,
		27129	=>	49632,
		27130	=>	49630,
		27131	=>	49627,
		27132	=>	49624,
		27133	=>	49621,
		27134	=>	49619,
		27135	=>	49616,
		27136	=>	49613,
		27137	=>	49611,
		27138	=>	49608,
		27139	=>	49605,
		27140	=>	49603,
		27141	=>	49600,
		27142	=>	49597,
		27143	=>	49594,
		27144	=>	49592,
		27145	=>	49589,
		27146	=>	49586,
		27147	=>	49584,
		27148	=>	49581,
		27149	=>	49578,
		27150	=>	49576,
		27151	=>	49573,
		27152	=>	49570,
		27153	=>	49568,
		27154	=>	49565,
		27155	=>	49562,
		27156	=>	49559,
		27157	=>	49557,
		27158	=>	49554,
		27159	=>	49551,
		27160	=>	49549,
		27161	=>	49546,
		27162	=>	49543,
		27163	=>	49541,
		27164	=>	49538,
		27165	=>	49535,
		27166	=>	49532,
		27167	=>	49530,
		27168	=>	49527,
		27169	=>	49524,
		27170	=>	49522,
		27171	=>	49519,
		27172	=>	49516,
		27173	=>	49514,
		27174	=>	49511,
		27175	=>	49508,
		27176	=>	49505,
		27177	=>	49503,
		27178	=>	49500,
		27179	=>	49497,
		27180	=>	49495,
		27181	=>	49492,
		27182	=>	49489,
		27183	=>	49487,
		27184	=>	49484,
		27185	=>	49481,
		27186	=>	49478,
		27187	=>	49476,
		27188	=>	49473,
		27189	=>	49470,
		27190	=>	49468,
		27191	=>	49465,
		27192	=>	49462,
		27193	=>	49460,
		27194	=>	49457,
		27195	=>	49454,
		27196	=>	49451,
		27197	=>	49449,
		27198	=>	49446,
		27199	=>	49443,
		27200	=>	49441,
		27201	=>	49438,
		27202	=>	49435,
		27203	=>	49432,
		27204	=>	49430,
		27205	=>	49427,
		27206	=>	49424,
		27207	=>	49422,
		27208	=>	49419,
		27209	=>	49416,
		27210	=>	49414,
		27211	=>	49411,
		27212	=>	49408,
		27213	=>	49405,
		27214	=>	49403,
		27215	=>	49400,
		27216	=>	49397,
		27217	=>	49395,
		27218	=>	49392,
		27219	=>	49389,
		27220	=>	49386,
		27221	=>	49384,
		27222	=>	49381,
		27223	=>	49378,
		27224	=>	49376,
		27225	=>	49373,
		27226	=>	49370,
		27227	=>	49368,
		27228	=>	49365,
		27229	=>	49362,
		27230	=>	49359,
		27231	=>	49357,
		27232	=>	49354,
		27233	=>	49351,
		27234	=>	49349,
		27235	=>	49346,
		27236	=>	49343,
		27237	=>	49340,
		27238	=>	49338,
		27239	=>	49335,
		27240	=>	49332,
		27241	=>	49330,
		27242	=>	49327,
		27243	=>	49324,
		27244	=>	49321,
		27245	=>	49319,
		27246	=>	49316,
		27247	=>	49313,
		27248	=>	49311,
		27249	=>	49308,
		27250	=>	49305,
		27251	=>	49302,
		27252	=>	49300,
		27253	=>	49297,
		27254	=>	49294,
		27255	=>	49292,
		27256	=>	49289,
		27257	=>	49286,
		27258	=>	49283,
		27259	=>	49281,
		27260	=>	49278,
		27261	=>	49275,
		27262	=>	49273,
		27263	=>	49270,
		27264	=>	49267,
		27265	=>	49264,
		27266	=>	49262,
		27267	=>	49259,
		27268	=>	49256,
		27269	=>	49254,
		27270	=>	49251,
		27271	=>	49248,
		27272	=>	49245,
		27273	=>	49243,
		27274	=>	49240,
		27275	=>	49237,
		27276	=>	49235,
		27277	=>	49232,
		27278	=>	49229,
		27279	=>	49226,
		27280	=>	49224,
		27281	=>	49221,
		27282	=>	49218,
		27283	=>	49216,
		27284	=>	49213,
		27285	=>	49210,
		27286	=>	49207,
		27287	=>	49205,
		27288	=>	49202,
		27289	=>	49199,
		27290	=>	49197,
		27291	=>	49194,
		27292	=>	49191,
		27293	=>	49188,
		27294	=>	49186,
		27295	=>	49183,
		27296	=>	49180,
		27297	=>	49178,
		27298	=>	49175,
		27299	=>	49172,
		27300	=>	49169,
		27301	=>	49167,
		27302	=>	49164,
		27303	=>	49161,
		27304	=>	49159,
		27305	=>	49156,
		27306	=>	49153,
		27307	=>	49150,
		27308	=>	49148,
		27309	=>	49145,
		27310	=>	49142,
		27311	=>	49139,
		27312	=>	49137,
		27313	=>	49134,
		27314	=>	49131,
		27315	=>	49129,
		27316	=>	49126,
		27317	=>	49123,
		27318	=>	49120,
		27319	=>	49118,
		27320	=>	49115,
		27321	=>	49112,
		27322	=>	49110,
		27323	=>	49107,
		27324	=>	49104,
		27325	=>	49101,
		27326	=>	49099,
		27327	=>	49096,
		27328	=>	49093,
		27329	=>	49090,
		27330	=>	49088,
		27331	=>	49085,
		27332	=>	49082,
		27333	=>	49080,
		27334	=>	49077,
		27335	=>	49074,
		27336	=>	49071,
		27337	=>	49069,
		27338	=>	49066,
		27339	=>	49063,
		27340	=>	49060,
		27341	=>	49058,
		27342	=>	49055,
		27343	=>	49052,
		27344	=>	49050,
		27345	=>	49047,
		27346	=>	49044,
		27347	=>	49041,
		27348	=>	49039,
		27349	=>	49036,
		27350	=>	49033,
		27351	=>	49030,
		27352	=>	49028,
		27353	=>	49025,
		27354	=>	49022,
		27355	=>	49020,
		27356	=>	49017,
		27357	=>	49014,
		27358	=>	49011,
		27359	=>	49009,
		27360	=>	49006,
		27361	=>	49003,
		27362	=>	49000,
		27363	=>	48998,
		27364	=>	48995,
		27365	=>	48992,
		27366	=>	48990,
		27367	=>	48987,
		27368	=>	48984,
		27369	=>	48981,
		27370	=>	48979,
		27371	=>	48976,
		27372	=>	48973,
		27373	=>	48970,
		27374	=>	48968,
		27375	=>	48965,
		27376	=>	48962,
		27377	=>	48960,
		27378	=>	48957,
		27379	=>	48954,
		27380	=>	48951,
		27381	=>	48949,
		27382	=>	48946,
		27383	=>	48943,
		27384	=>	48940,
		27385	=>	48938,
		27386	=>	48935,
		27387	=>	48932,
		27388	=>	48929,
		27389	=>	48927,
		27390	=>	48924,
		27391	=>	48921,
		27392	=>	48919,
		27393	=>	48916,
		27394	=>	48913,
		27395	=>	48910,
		27396	=>	48908,
		27397	=>	48905,
		27398	=>	48902,
		27399	=>	48899,
		27400	=>	48897,
		27401	=>	48894,
		27402	=>	48891,
		27403	=>	48888,
		27404	=>	48886,
		27405	=>	48883,
		27406	=>	48880,
		27407	=>	48878,
		27408	=>	48875,
		27409	=>	48872,
		27410	=>	48869,
		27411	=>	48867,
		27412	=>	48864,
		27413	=>	48861,
		27414	=>	48858,
		27415	=>	48856,
		27416	=>	48853,
		27417	=>	48850,
		27418	=>	48847,
		27419	=>	48845,
		27420	=>	48842,
		27421	=>	48839,
		27422	=>	48836,
		27423	=>	48834,
		27424	=>	48831,
		27425	=>	48828,
		27426	=>	48826,
		27427	=>	48823,
		27428	=>	48820,
		27429	=>	48817,
		27430	=>	48815,
		27431	=>	48812,
		27432	=>	48809,
		27433	=>	48806,
		27434	=>	48804,
		27435	=>	48801,
		27436	=>	48798,
		27437	=>	48795,
		27438	=>	48793,
		27439	=>	48790,
		27440	=>	48787,
		27441	=>	48784,
		27442	=>	48782,
		27443	=>	48779,
		27444	=>	48776,
		27445	=>	48773,
		27446	=>	48771,
		27447	=>	48768,
		27448	=>	48765,
		27449	=>	48762,
		27450	=>	48760,
		27451	=>	48757,
		27452	=>	48754,
		27453	=>	48752,
		27454	=>	48749,
		27455	=>	48746,
		27456	=>	48743,
		27457	=>	48741,
		27458	=>	48738,
		27459	=>	48735,
		27460	=>	48732,
		27461	=>	48730,
		27462	=>	48727,
		27463	=>	48724,
		27464	=>	48721,
		27465	=>	48719,
		27466	=>	48716,
		27467	=>	48713,
		27468	=>	48710,
		27469	=>	48708,
		27470	=>	48705,
		27471	=>	48702,
		27472	=>	48699,
		27473	=>	48697,
		27474	=>	48694,
		27475	=>	48691,
		27476	=>	48688,
		27477	=>	48686,
		27478	=>	48683,
		27479	=>	48680,
		27480	=>	48677,
		27481	=>	48675,
		27482	=>	48672,
		27483	=>	48669,
		27484	=>	48666,
		27485	=>	48664,
		27486	=>	48661,
		27487	=>	48658,
		27488	=>	48655,
		27489	=>	48653,
		27490	=>	48650,
		27491	=>	48647,
		27492	=>	48644,
		27493	=>	48642,
		27494	=>	48639,
		27495	=>	48636,
		27496	=>	48633,
		27497	=>	48631,
		27498	=>	48628,
		27499	=>	48625,
		27500	=>	48622,
		27501	=>	48620,
		27502	=>	48617,
		27503	=>	48614,
		27504	=>	48611,
		27505	=>	48609,
		27506	=>	48606,
		27507	=>	48603,
		27508	=>	48600,
		27509	=>	48598,
		27510	=>	48595,
		27511	=>	48592,
		27512	=>	48589,
		27513	=>	48587,
		27514	=>	48584,
		27515	=>	48581,
		27516	=>	48578,
		27517	=>	48576,
		27518	=>	48573,
		27519	=>	48570,
		27520	=>	48567,
		27521	=>	48565,
		27522	=>	48562,
		27523	=>	48559,
		27524	=>	48556,
		27525	=>	48554,
		27526	=>	48551,
		27527	=>	48548,
		27528	=>	48545,
		27529	=>	48543,
		27530	=>	48540,
		27531	=>	48537,
		27532	=>	48534,
		27533	=>	48532,
		27534	=>	48529,
		27535	=>	48526,
		27536	=>	48523,
		27537	=>	48521,
		27538	=>	48518,
		27539	=>	48515,
		27540	=>	48512,
		27541	=>	48510,
		27542	=>	48507,
		27543	=>	48504,
		27544	=>	48501,
		27545	=>	48499,
		27546	=>	48496,
		27547	=>	48493,
		27548	=>	48490,
		27549	=>	48488,
		27550	=>	48485,
		27551	=>	48482,
		27552	=>	48479,
		27553	=>	48477,
		27554	=>	48474,
		27555	=>	48471,
		27556	=>	48468,
		27557	=>	48466,
		27558	=>	48463,
		27559	=>	48460,
		27560	=>	48457,
		27561	=>	48454,
		27562	=>	48452,
		27563	=>	48449,
		27564	=>	48446,
		27565	=>	48443,
		27566	=>	48441,
		27567	=>	48438,
		27568	=>	48435,
		27569	=>	48432,
		27570	=>	48430,
		27571	=>	48427,
		27572	=>	48424,
		27573	=>	48421,
		27574	=>	48419,
		27575	=>	48416,
		27576	=>	48413,
		27577	=>	48410,
		27578	=>	48408,
		27579	=>	48405,
		27580	=>	48402,
		27581	=>	48399,
		27582	=>	48397,
		27583	=>	48394,
		27584	=>	48391,
		27585	=>	48388,
		27586	=>	48385,
		27587	=>	48383,
		27588	=>	48380,
		27589	=>	48377,
		27590	=>	48374,
		27591	=>	48372,
		27592	=>	48369,
		27593	=>	48366,
		27594	=>	48363,
		27595	=>	48361,
		27596	=>	48358,
		27597	=>	48355,
		27598	=>	48352,
		27599	=>	48350,
		27600	=>	48347,
		27601	=>	48344,
		27602	=>	48341,
		27603	=>	48339,
		27604	=>	48336,
		27605	=>	48333,
		27606	=>	48330,
		27607	=>	48327,
		27608	=>	48325,
		27609	=>	48322,
		27610	=>	48319,
		27611	=>	48316,
		27612	=>	48314,
		27613	=>	48311,
		27614	=>	48308,
		27615	=>	48305,
		27616	=>	48303,
		27617	=>	48300,
		27618	=>	48297,
		27619	=>	48294,
		27620	=>	48292,
		27621	=>	48289,
		27622	=>	48286,
		27623	=>	48283,
		27624	=>	48280,
		27625	=>	48278,
		27626	=>	48275,
		27627	=>	48272,
		27628	=>	48269,
		27629	=>	48267,
		27630	=>	48264,
		27631	=>	48261,
		27632	=>	48258,
		27633	=>	48256,
		27634	=>	48253,
		27635	=>	48250,
		27636	=>	48247,
		27637	=>	48244,
		27638	=>	48242,
		27639	=>	48239,
		27640	=>	48236,
		27641	=>	48233,
		27642	=>	48231,
		27643	=>	48228,
		27644	=>	48225,
		27645	=>	48222,
		27646	=>	48220,
		27647	=>	48217,
		27648	=>	48214,
		27649	=>	48211,
		27650	=>	48208,
		27651	=>	48206,
		27652	=>	48203,
		27653	=>	48200,
		27654	=>	48197,
		27655	=>	48195,
		27656	=>	48192,
		27657	=>	48189,
		27658	=>	48186,
		27659	=>	48184,
		27660	=>	48181,
		27661	=>	48178,
		27662	=>	48175,
		27663	=>	48172,
		27664	=>	48170,
		27665	=>	48167,
		27666	=>	48164,
		27667	=>	48161,
		27668	=>	48159,
		27669	=>	48156,
		27670	=>	48153,
		27671	=>	48150,
		27672	=>	48147,
		27673	=>	48145,
		27674	=>	48142,
		27675	=>	48139,
		27676	=>	48136,
		27677	=>	48134,
		27678	=>	48131,
		27679	=>	48128,
		27680	=>	48125,
		27681	=>	48122,
		27682	=>	48120,
		27683	=>	48117,
		27684	=>	48114,
		27685	=>	48111,
		27686	=>	48109,
		27687	=>	48106,
		27688	=>	48103,
		27689	=>	48100,
		27690	=>	48098,
		27691	=>	48095,
		27692	=>	48092,
		27693	=>	48089,
		27694	=>	48086,
		27695	=>	48084,
		27696	=>	48081,
		27697	=>	48078,
		27698	=>	48075,
		27699	=>	48073,
		27700	=>	48070,
		27701	=>	48067,
		27702	=>	48064,
		27703	=>	48061,
		27704	=>	48059,
		27705	=>	48056,
		27706	=>	48053,
		27707	=>	48050,
		27708	=>	48048,
		27709	=>	48045,
		27710	=>	48042,
		27711	=>	48039,
		27712	=>	48036,
		27713	=>	48034,
		27714	=>	48031,
		27715	=>	48028,
		27716	=>	48025,
		27717	=>	48022,
		27718	=>	48020,
		27719	=>	48017,
		27720	=>	48014,
		27721	=>	48011,
		27722	=>	48009,
		27723	=>	48006,
		27724	=>	48003,
		27725	=>	48000,
		27726	=>	47997,
		27727	=>	47995,
		27728	=>	47992,
		27729	=>	47989,
		27730	=>	47986,
		27731	=>	47984,
		27732	=>	47981,
		27733	=>	47978,
		27734	=>	47975,
		27735	=>	47972,
		27736	=>	47970,
		27737	=>	47967,
		27738	=>	47964,
		27739	=>	47961,
		27740	=>	47959,
		27741	=>	47956,
		27742	=>	47953,
		27743	=>	47950,
		27744	=>	47947,
		27745	=>	47945,
		27746	=>	47942,
		27747	=>	47939,
		27748	=>	47936,
		27749	=>	47933,
		27750	=>	47931,
		27751	=>	47928,
		27752	=>	47925,
		27753	=>	47922,
		27754	=>	47920,
		27755	=>	47917,
		27756	=>	47914,
		27757	=>	47911,
		27758	=>	47908,
		27759	=>	47906,
		27760	=>	47903,
		27761	=>	47900,
		27762	=>	47897,
		27763	=>	47894,
		27764	=>	47892,
		27765	=>	47889,
		27766	=>	47886,
		27767	=>	47883,
		27768	=>	47881,
		27769	=>	47878,
		27770	=>	47875,
		27771	=>	47872,
		27772	=>	47869,
		27773	=>	47867,
		27774	=>	47864,
		27775	=>	47861,
		27776	=>	47858,
		27777	=>	47855,
		27778	=>	47853,
		27779	=>	47850,
		27780	=>	47847,
		27781	=>	47844,
		27782	=>	47841,
		27783	=>	47839,
		27784	=>	47836,
		27785	=>	47833,
		27786	=>	47830,
		27787	=>	47828,
		27788	=>	47825,
		27789	=>	47822,
		27790	=>	47819,
		27791	=>	47816,
		27792	=>	47814,
		27793	=>	47811,
		27794	=>	47808,
		27795	=>	47805,
		27796	=>	47802,
		27797	=>	47800,
		27798	=>	47797,
		27799	=>	47794,
		27800	=>	47791,
		27801	=>	47788,
		27802	=>	47786,
		27803	=>	47783,
		27804	=>	47780,
		27805	=>	47777,
		27806	=>	47774,
		27807	=>	47772,
		27808	=>	47769,
		27809	=>	47766,
		27810	=>	47763,
		27811	=>	47761,
		27812	=>	47758,
		27813	=>	47755,
		27814	=>	47752,
		27815	=>	47749,
		27816	=>	47747,
		27817	=>	47744,
		27818	=>	47741,
		27819	=>	47738,
		27820	=>	47735,
		27821	=>	47733,
		27822	=>	47730,
		27823	=>	47727,
		27824	=>	47724,
		27825	=>	47721,
		27826	=>	47719,
		27827	=>	47716,
		27828	=>	47713,
		27829	=>	47710,
		27830	=>	47707,
		27831	=>	47705,
		27832	=>	47702,
		27833	=>	47699,
		27834	=>	47696,
		27835	=>	47693,
		27836	=>	47691,
		27837	=>	47688,
		27838	=>	47685,
		27839	=>	47682,
		27840	=>	47679,
		27841	=>	47677,
		27842	=>	47674,
		27843	=>	47671,
		27844	=>	47668,
		27845	=>	47665,
		27846	=>	47663,
		27847	=>	47660,
		27848	=>	47657,
		27849	=>	47654,
		27850	=>	47651,
		27851	=>	47649,
		27852	=>	47646,
		27853	=>	47643,
		27854	=>	47640,
		27855	=>	47637,
		27856	=>	47635,
		27857	=>	47632,
		27858	=>	47629,
		27859	=>	47626,
		27860	=>	47623,
		27861	=>	47621,
		27862	=>	47618,
		27863	=>	47615,
		27864	=>	47612,
		27865	=>	47609,
		27866	=>	47607,
		27867	=>	47604,
		27868	=>	47601,
		27869	=>	47598,
		27870	=>	47595,
		27871	=>	47593,
		27872	=>	47590,
		27873	=>	47587,
		27874	=>	47584,
		27875	=>	47581,
		27876	=>	47579,
		27877	=>	47576,
		27878	=>	47573,
		27879	=>	47570,
		27880	=>	47567,
		27881	=>	47565,
		27882	=>	47562,
		27883	=>	47559,
		27884	=>	47556,
		27885	=>	47553,
		27886	=>	47551,
		27887	=>	47548,
		27888	=>	47545,
		27889	=>	47542,
		27890	=>	47539,
		27891	=>	47537,
		27892	=>	47534,
		27893	=>	47531,
		27894	=>	47528,
		27895	=>	47525,
		27896	=>	47523,
		27897	=>	47520,
		27898	=>	47517,
		27899	=>	47514,
		27900	=>	47511,
		27901	=>	47509,
		27902	=>	47506,
		27903	=>	47503,
		27904	=>	47500,
		27905	=>	47497,
		27906	=>	47495,
		27907	=>	47492,
		27908	=>	47489,
		27909	=>	47486,
		27910	=>	47483,
		27911	=>	47480,
		27912	=>	47478,
		27913	=>	47475,
		27914	=>	47472,
		27915	=>	47469,
		27916	=>	47466,
		27917	=>	47464,
		27918	=>	47461,
		27919	=>	47458,
		27920	=>	47455,
		27921	=>	47452,
		27922	=>	47450,
		27923	=>	47447,
		27924	=>	47444,
		27925	=>	47441,
		27926	=>	47438,
		27927	=>	47436,
		27928	=>	47433,
		27929	=>	47430,
		27930	=>	47427,
		27931	=>	47424,
		27932	=>	47422,
		27933	=>	47419,
		27934	=>	47416,
		27935	=>	47413,
		27936	=>	47410,
		27937	=>	47407,
		27938	=>	47405,
		27939	=>	47402,
		27940	=>	47399,
		27941	=>	47396,
		27942	=>	47393,
		27943	=>	47391,
		27944	=>	47388,
		27945	=>	47385,
		27946	=>	47382,
		27947	=>	47379,
		27948	=>	47377,
		27949	=>	47374,
		27950	=>	47371,
		27951	=>	47368,
		27952	=>	47365,
		27953	=>	47362,
		27954	=>	47360,
		27955	=>	47357,
		27956	=>	47354,
		27957	=>	47351,
		27958	=>	47348,
		27959	=>	47346,
		27960	=>	47343,
		27961	=>	47340,
		27962	=>	47337,
		27963	=>	47334,
		27964	=>	47332,
		27965	=>	47329,
		27966	=>	47326,
		27967	=>	47323,
		27968	=>	47320,
		27969	=>	47317,
		27970	=>	47315,
		27971	=>	47312,
		27972	=>	47309,
		27973	=>	47306,
		27974	=>	47303,
		27975	=>	47301,
		27976	=>	47298,
		27977	=>	47295,
		27978	=>	47292,
		27979	=>	47289,
		27980	=>	47286,
		27981	=>	47284,
		27982	=>	47281,
		27983	=>	47278,
		27984	=>	47275,
		27985	=>	47272,
		27986	=>	47270,
		27987	=>	47267,
		27988	=>	47264,
		27989	=>	47261,
		27990	=>	47258,
		27991	=>	47255,
		27992	=>	47253,
		27993	=>	47250,
		27994	=>	47247,
		27995	=>	47244,
		27996	=>	47241,
		27997	=>	47239,
		27998	=>	47236,
		27999	=>	47233,
		28000	=>	47230,
		28001	=>	47227,
		28002	=>	47224,
		28003	=>	47222,
		28004	=>	47219,
		28005	=>	47216,
		28006	=>	47213,
		28007	=>	47210,
		28008	=>	47208,
		28009	=>	47205,
		28010	=>	47202,
		28011	=>	47199,
		28012	=>	47196,
		28013	=>	47193,
		28014	=>	47191,
		28015	=>	47188,
		28016	=>	47185,
		28017	=>	47182,
		28018	=>	47179,
		28019	=>	47177,
		28020	=>	47174,
		28021	=>	47171,
		28022	=>	47168,
		28023	=>	47165,
		28024	=>	47162,
		28025	=>	47160,
		28026	=>	47157,
		28027	=>	47154,
		28028	=>	47151,
		28029	=>	47148,
		28030	=>	47146,
		28031	=>	47143,
		28032	=>	47140,
		28033	=>	47137,
		28034	=>	47134,
		28035	=>	47131,
		28036	=>	47129,
		28037	=>	47126,
		28038	=>	47123,
		28039	=>	47120,
		28040	=>	47117,
		28041	=>	47114,
		28042	=>	47112,
		28043	=>	47109,
		28044	=>	47106,
		28045	=>	47103,
		28046	=>	47100,
		28047	=>	47097,
		28048	=>	47095,
		28049	=>	47092,
		28050	=>	47089,
		28051	=>	47086,
		28052	=>	47083,
		28053	=>	47081,
		28054	=>	47078,
		28055	=>	47075,
		28056	=>	47072,
		28057	=>	47069,
		28058	=>	47066,
		28059	=>	47064,
		28060	=>	47061,
		28061	=>	47058,
		28062	=>	47055,
		28063	=>	47052,
		28064	=>	47049,
		28065	=>	47047,
		28066	=>	47044,
		28067	=>	47041,
		28068	=>	47038,
		28069	=>	47035,
		28070	=>	47032,
		28071	=>	47030,
		28072	=>	47027,
		28073	=>	47024,
		28074	=>	47021,
		28075	=>	47018,
		28076	=>	47016,
		28077	=>	47013,
		28078	=>	47010,
		28079	=>	47007,
		28080	=>	47004,
		28081	=>	47001,
		28082	=>	46999,
		28083	=>	46996,
		28084	=>	46993,
		28085	=>	46990,
		28086	=>	46987,
		28087	=>	46984,
		28088	=>	46982,
		28089	=>	46979,
		28090	=>	46976,
		28091	=>	46973,
		28092	=>	46970,
		28093	=>	46967,
		28094	=>	46965,
		28095	=>	46962,
		28096	=>	46959,
		28097	=>	46956,
		28098	=>	46953,
		28099	=>	46950,
		28100	=>	46948,
		28101	=>	46945,
		28102	=>	46942,
		28103	=>	46939,
		28104	=>	46936,
		28105	=>	46933,
		28106	=>	46931,
		28107	=>	46928,
		28108	=>	46925,
		28109	=>	46922,
		28110	=>	46919,
		28111	=>	46916,
		28112	=>	46914,
		28113	=>	46911,
		28114	=>	46908,
		28115	=>	46905,
		28116	=>	46902,
		28117	=>	46899,
		28118	=>	46897,
		28119	=>	46894,
		28120	=>	46891,
		28121	=>	46888,
		28122	=>	46885,
		28123	=>	46882,
		28124	=>	46880,
		28125	=>	46877,
		28126	=>	46874,
		28127	=>	46871,
		28128	=>	46868,
		28129	=>	46865,
		28130	=>	46863,
		28131	=>	46860,
		28132	=>	46857,
		28133	=>	46854,
		28134	=>	46851,
		28135	=>	46848,
		28136	=>	46846,
		28137	=>	46843,
		28138	=>	46840,
		28139	=>	46837,
		28140	=>	46834,
		28141	=>	46831,
		28142	=>	46829,
		28143	=>	46826,
		28144	=>	46823,
		28145	=>	46820,
		28146	=>	46817,
		28147	=>	46814,
		28148	=>	46811,
		28149	=>	46809,
		28150	=>	46806,
		28151	=>	46803,
		28152	=>	46800,
		28153	=>	46797,
		28154	=>	46794,
		28155	=>	46792,
		28156	=>	46789,
		28157	=>	46786,
		28158	=>	46783,
		28159	=>	46780,
		28160	=>	46777,
		28161	=>	46775,
		28162	=>	46772,
		28163	=>	46769,
		28164	=>	46766,
		28165	=>	46763,
		28166	=>	46760,
		28167	=>	46758,
		28168	=>	46755,
		28169	=>	46752,
		28170	=>	46749,
		28171	=>	46746,
		28172	=>	46743,
		28173	=>	46740,
		28174	=>	46738,
		28175	=>	46735,
		28176	=>	46732,
		28177	=>	46729,
		28178	=>	46726,
		28179	=>	46723,
		28180	=>	46721,
		28181	=>	46718,
		28182	=>	46715,
		28183	=>	46712,
		28184	=>	46709,
		28185	=>	46706,
		28186	=>	46704,
		28187	=>	46701,
		28188	=>	46698,
		28189	=>	46695,
		28190	=>	46692,
		28191	=>	46689,
		28192	=>	46686,
		28193	=>	46684,
		28194	=>	46681,
		28195	=>	46678,
		28196	=>	46675,
		28197	=>	46672,
		28198	=>	46669,
		28199	=>	46667,
		28200	=>	46664,
		28201	=>	46661,
		28202	=>	46658,
		28203	=>	46655,
		28204	=>	46652,
		28205	=>	46649,
		28206	=>	46647,
		28207	=>	46644,
		28208	=>	46641,
		28209	=>	46638,
		28210	=>	46635,
		28211	=>	46632,
		28212	=>	46630,
		28213	=>	46627,
		28214	=>	46624,
		28215	=>	46621,
		28216	=>	46618,
		28217	=>	46615,
		28218	=>	46612,
		28219	=>	46610,
		28220	=>	46607,
		28221	=>	46604,
		28222	=>	46601,
		28223	=>	46598,
		28224	=>	46595,
		28225	=>	46593,
		28226	=>	46590,
		28227	=>	46587,
		28228	=>	46584,
		28229	=>	46581,
		28230	=>	46578,
		28231	=>	46575,
		28232	=>	46573,
		28233	=>	46570,
		28234	=>	46567,
		28235	=>	46564,
		28236	=>	46561,
		28237	=>	46558,
		28238	=>	46556,
		28239	=>	46553,
		28240	=>	46550,
		28241	=>	46547,
		28242	=>	46544,
		28243	=>	46541,
		28244	=>	46538,
		28245	=>	46536,
		28246	=>	46533,
		28247	=>	46530,
		28248	=>	46527,
		28249	=>	46524,
		28250	=>	46521,
		28251	=>	46518,
		28252	=>	46516,
		28253	=>	46513,
		28254	=>	46510,
		28255	=>	46507,
		28256	=>	46504,
		28257	=>	46501,
		28258	=>	46498,
		28259	=>	46496,
		28260	=>	46493,
		28261	=>	46490,
		28262	=>	46487,
		28263	=>	46484,
		28264	=>	46481,
		28265	=>	46479,
		28266	=>	46476,
		28267	=>	46473,
		28268	=>	46470,
		28269	=>	46467,
		28270	=>	46464,
		28271	=>	46461,
		28272	=>	46459,
		28273	=>	46456,
		28274	=>	46453,
		28275	=>	46450,
		28276	=>	46447,
		28277	=>	46444,
		28278	=>	46441,
		28279	=>	46439,
		28280	=>	46436,
		28281	=>	46433,
		28282	=>	46430,
		28283	=>	46427,
		28284	=>	46424,
		28285	=>	46421,
		28286	=>	46419,
		28287	=>	46416,
		28288	=>	46413,
		28289	=>	46410,
		28290	=>	46407,
		28291	=>	46404,
		28292	=>	46401,
		28293	=>	46399,
		28294	=>	46396,
		28295	=>	46393,
		28296	=>	46390,
		28297	=>	46387,
		28298	=>	46384,
		28299	=>	46381,
		28300	=>	46379,
		28301	=>	46376,
		28302	=>	46373,
		28303	=>	46370,
		28304	=>	46367,
		28305	=>	46364,
		28306	=>	46361,
		28307	=>	46359,
		28308	=>	46356,
		28309	=>	46353,
		28310	=>	46350,
		28311	=>	46347,
		28312	=>	46344,
		28313	=>	46341,
		28314	=>	46339,
		28315	=>	46336,
		28316	=>	46333,
		28317	=>	46330,
		28318	=>	46327,
		28319	=>	46324,
		28320	=>	46321,
		28321	=>	46319,
		28322	=>	46316,
		28323	=>	46313,
		28324	=>	46310,
		28325	=>	46307,
		28326	=>	46304,
		28327	=>	46301,
		28328	=>	46299,
		28329	=>	46296,
		28330	=>	46293,
		28331	=>	46290,
		28332	=>	46287,
		28333	=>	46284,
		28334	=>	46281,
		28335	=>	46278,
		28336	=>	46276,
		28337	=>	46273,
		28338	=>	46270,
		28339	=>	46267,
		28340	=>	46264,
		28341	=>	46261,
		28342	=>	46258,
		28343	=>	46256,
		28344	=>	46253,
		28345	=>	46250,
		28346	=>	46247,
		28347	=>	46244,
		28348	=>	46241,
		28349	=>	46238,
		28350	=>	46236,
		28351	=>	46233,
		28352	=>	46230,
		28353	=>	46227,
		28354	=>	46224,
		28355	=>	46221,
		28356	=>	46218,
		28357	=>	46215,
		28358	=>	46213,
		28359	=>	46210,
		28360	=>	46207,
		28361	=>	46204,
		28362	=>	46201,
		28363	=>	46198,
		28364	=>	46195,
		28365	=>	46193,
		28366	=>	46190,
		28367	=>	46187,
		28368	=>	46184,
		28369	=>	46181,
		28370	=>	46178,
		28371	=>	46175,
		28372	=>	46172,
		28373	=>	46170,
		28374	=>	46167,
		28375	=>	46164,
		28376	=>	46161,
		28377	=>	46158,
		28378	=>	46155,
		28379	=>	46152,
		28380	=>	46150,
		28381	=>	46147,
		28382	=>	46144,
		28383	=>	46141,
		28384	=>	46138,
		28385	=>	46135,
		28386	=>	46132,
		28387	=>	46129,
		28388	=>	46127,
		28389	=>	46124,
		28390	=>	46121,
		28391	=>	46118,
		28392	=>	46115,
		28393	=>	46112,
		28394	=>	46109,
		28395	=>	46107,
		28396	=>	46104,
		28397	=>	46101,
		28398	=>	46098,
		28399	=>	46095,
		28400	=>	46092,
		28401	=>	46089,
		28402	=>	46086,
		28403	=>	46084,
		28404	=>	46081,
		28405	=>	46078,
		28406	=>	46075,
		28407	=>	46072,
		28408	=>	46069,
		28409	=>	46066,
		28410	=>	46063,
		28411	=>	46061,
		28412	=>	46058,
		28413	=>	46055,
		28414	=>	46052,
		28415	=>	46049,
		28416	=>	46046,
		28417	=>	46043,
		28418	=>	46041,
		28419	=>	46038,
		28420	=>	46035,
		28421	=>	46032,
		28422	=>	46029,
		28423	=>	46026,
		28424	=>	46023,
		28425	=>	46020,
		28426	=>	46018,
		28427	=>	46015,
		28428	=>	46012,
		28429	=>	46009,
		28430	=>	46006,
		28431	=>	46003,
		28432	=>	46000,
		28433	=>	45997,
		28434	=>	45995,
		28435	=>	45992,
		28436	=>	45989,
		28437	=>	45986,
		28438	=>	45983,
		28439	=>	45980,
		28440	=>	45977,
		28441	=>	45974,
		28442	=>	45972,
		28443	=>	45969,
		28444	=>	45966,
		28445	=>	45963,
		28446	=>	45960,
		28447	=>	45957,
		28448	=>	45954,
		28449	=>	45951,
		28450	=>	45949,
		28451	=>	45946,
		28452	=>	45943,
		28453	=>	45940,
		28454	=>	45937,
		28455	=>	45934,
		28456	=>	45931,
		28457	=>	45928,
		28458	=>	45926,
		28459	=>	45923,
		28460	=>	45920,
		28461	=>	45917,
		28462	=>	45914,
		28463	=>	45911,
		28464	=>	45908,
		28465	=>	45905,
		28466	=>	45902,
		28467	=>	45900,
		28468	=>	45897,
		28469	=>	45894,
		28470	=>	45891,
		28471	=>	45888,
		28472	=>	45885,
		28473	=>	45882,
		28474	=>	45879,
		28475	=>	45877,
		28476	=>	45874,
		28477	=>	45871,
		28478	=>	45868,
		28479	=>	45865,
		28480	=>	45862,
		28481	=>	45859,
		28482	=>	45856,
		28483	=>	45854,
		28484	=>	45851,
		28485	=>	45848,
		28486	=>	45845,
		28487	=>	45842,
		28488	=>	45839,
		28489	=>	45836,
		28490	=>	45833,
		28491	=>	45831,
		28492	=>	45828,
		28493	=>	45825,
		28494	=>	45822,
		28495	=>	45819,
		28496	=>	45816,
		28497	=>	45813,
		28498	=>	45810,
		28499	=>	45807,
		28500	=>	45805,
		28501	=>	45802,
		28502	=>	45799,
		28503	=>	45796,
		28504	=>	45793,
		28505	=>	45790,
		28506	=>	45787,
		28507	=>	45784,
		28508	=>	45782,
		28509	=>	45779,
		28510	=>	45776,
		28511	=>	45773,
		28512	=>	45770,
		28513	=>	45767,
		28514	=>	45764,
		28515	=>	45761,
		28516	=>	45758,
		28517	=>	45756,
		28518	=>	45753,
		28519	=>	45750,
		28520	=>	45747,
		28521	=>	45744,
		28522	=>	45741,
		28523	=>	45738,
		28524	=>	45735,
		28525	=>	45732,
		28526	=>	45730,
		28527	=>	45727,
		28528	=>	45724,
		28529	=>	45721,
		28530	=>	45718,
		28531	=>	45715,
		28532	=>	45712,
		28533	=>	45709,
		28534	=>	45707,
		28535	=>	45704,
		28536	=>	45701,
		28537	=>	45698,
		28538	=>	45695,
		28539	=>	45692,
		28540	=>	45689,
		28541	=>	45686,
		28542	=>	45683,
		28543	=>	45681,
		28544	=>	45678,
		28545	=>	45675,
		28546	=>	45672,
		28547	=>	45669,
		28548	=>	45666,
		28549	=>	45663,
		28550	=>	45660,
		28551	=>	45657,
		28552	=>	45655,
		28553	=>	45652,
		28554	=>	45649,
		28555	=>	45646,
		28556	=>	45643,
		28557	=>	45640,
		28558	=>	45637,
		28559	=>	45634,
		28560	=>	45631,
		28561	=>	45629,
		28562	=>	45626,
		28563	=>	45623,
		28564	=>	45620,
		28565	=>	45617,
		28566	=>	45614,
		28567	=>	45611,
		28568	=>	45608,
		28569	=>	45605,
		28570	=>	45603,
		28571	=>	45600,
		28572	=>	45597,
		28573	=>	45594,
		28574	=>	45591,
		28575	=>	45588,
		28576	=>	45585,
		28577	=>	45582,
		28578	=>	45579,
		28579	=>	45577,
		28580	=>	45574,
		28581	=>	45571,
		28582	=>	45568,
		28583	=>	45565,
		28584	=>	45562,
		28585	=>	45559,
		28586	=>	45556,
		28587	=>	45553,
		28588	=>	45550,
		28589	=>	45548,
		28590	=>	45545,
		28591	=>	45542,
		28592	=>	45539,
		28593	=>	45536,
		28594	=>	45533,
		28595	=>	45530,
		28596	=>	45527,
		28597	=>	45524,
		28598	=>	45522,
		28599	=>	45519,
		28600	=>	45516,
		28601	=>	45513,
		28602	=>	45510,
		28603	=>	45507,
		28604	=>	45504,
		28605	=>	45501,
		28606	=>	45498,
		28607	=>	45495,
		28608	=>	45493,
		28609	=>	45490,
		28610	=>	45487,
		28611	=>	45484,
		28612	=>	45481,
		28613	=>	45478,
		28614	=>	45475,
		28615	=>	45472,
		28616	=>	45469,
		28617	=>	45467,
		28618	=>	45464,
		28619	=>	45461,
		28620	=>	45458,
		28621	=>	45455,
		28622	=>	45452,
		28623	=>	45449,
		28624	=>	45446,
		28625	=>	45443,
		28626	=>	45440,
		28627	=>	45438,
		28628	=>	45435,
		28629	=>	45432,
		28630	=>	45429,
		28631	=>	45426,
		28632	=>	45423,
		28633	=>	45420,
		28634	=>	45417,
		28635	=>	45414,
		28636	=>	45411,
		28637	=>	45409,
		28638	=>	45406,
		28639	=>	45403,
		28640	=>	45400,
		28641	=>	45397,
		28642	=>	45394,
		28643	=>	45391,
		28644	=>	45388,
		28645	=>	45385,
		28646	=>	45383,
		28647	=>	45380,
		28648	=>	45377,
		28649	=>	45374,
		28650	=>	45371,
		28651	=>	45368,
		28652	=>	45365,
		28653	=>	45362,
		28654	=>	45359,
		28655	=>	45356,
		28656	=>	45354,
		28657	=>	45351,
		28658	=>	45348,
		28659	=>	45345,
		28660	=>	45342,
		28661	=>	45339,
		28662	=>	45336,
		28663	=>	45333,
		28664	=>	45330,
		28665	=>	45327,
		28666	=>	45324,
		28667	=>	45322,
		28668	=>	45319,
		28669	=>	45316,
		28670	=>	45313,
		28671	=>	45310,
		28672	=>	45307,
		28673	=>	45304,
		28674	=>	45301,
		28675	=>	45298,
		28676	=>	45295,
		28677	=>	45293,
		28678	=>	45290,
		28679	=>	45287,
		28680	=>	45284,
		28681	=>	45281,
		28682	=>	45278,
		28683	=>	45275,
		28684	=>	45272,
		28685	=>	45269,
		28686	=>	45266,
		28687	=>	45264,
		28688	=>	45261,
		28689	=>	45258,
		28690	=>	45255,
		28691	=>	45252,
		28692	=>	45249,
		28693	=>	45246,
		28694	=>	45243,
		28695	=>	45240,
		28696	=>	45237,
		28697	=>	45234,
		28698	=>	45232,
		28699	=>	45229,
		28700	=>	45226,
		28701	=>	45223,
		28702	=>	45220,
		28703	=>	45217,
		28704	=>	45214,
		28705	=>	45211,
		28706	=>	45208,
		28707	=>	45205,
		28708	=>	45203,
		28709	=>	45200,
		28710	=>	45197,
		28711	=>	45194,
		28712	=>	45191,
		28713	=>	45188,
		28714	=>	45185,
		28715	=>	45182,
		28716	=>	45179,
		28717	=>	45176,
		28718	=>	45173,
		28719	=>	45171,
		28720	=>	45168,
		28721	=>	45165,
		28722	=>	45162,
		28723	=>	45159,
		28724	=>	45156,
		28725	=>	45153,
		28726	=>	45150,
		28727	=>	45147,
		28728	=>	45144,
		28729	=>	45141,
		28730	=>	45139,
		28731	=>	45136,
		28732	=>	45133,
		28733	=>	45130,
		28734	=>	45127,
		28735	=>	45124,
		28736	=>	45121,
		28737	=>	45118,
		28738	=>	45115,
		28739	=>	45112,
		28740	=>	45109,
		28741	=>	45107,
		28742	=>	45104,
		28743	=>	45101,
		28744	=>	45098,
		28745	=>	45095,
		28746	=>	45092,
		28747	=>	45089,
		28748	=>	45086,
		28749	=>	45083,
		28750	=>	45080,
		28751	=>	45077,
		28752	=>	45075,
		28753	=>	45072,
		28754	=>	45069,
		28755	=>	45066,
		28756	=>	45063,
		28757	=>	45060,
		28758	=>	45057,
		28759	=>	45054,
		28760	=>	45051,
		28761	=>	45048,
		28762	=>	45045,
		28763	=>	45042,
		28764	=>	45040,
		28765	=>	45037,
		28766	=>	45034,
		28767	=>	45031,
		28768	=>	45028,
		28769	=>	45025,
		28770	=>	45022,
		28771	=>	45019,
		28772	=>	45016,
		28773	=>	45013,
		28774	=>	45010,
		28775	=>	45008,
		28776	=>	45005,
		28777	=>	45002,
		28778	=>	44999,
		28779	=>	44996,
		28780	=>	44993,
		28781	=>	44990,
		28782	=>	44987,
		28783	=>	44984,
		28784	=>	44981,
		28785	=>	44978,
		28786	=>	44975,
		28787	=>	44973,
		28788	=>	44970,
		28789	=>	44967,
		28790	=>	44964,
		28791	=>	44961,
		28792	=>	44958,
		28793	=>	44955,
		28794	=>	44952,
		28795	=>	44949,
		28796	=>	44946,
		28797	=>	44943,
		28798	=>	44940,
		28799	=>	44938,
		28800	=>	44935,
		28801	=>	44932,
		28802	=>	44929,
		28803	=>	44926,
		28804	=>	44923,
		28805	=>	44920,
		28806	=>	44917,
		28807	=>	44914,
		28808	=>	44911,
		28809	=>	44908,
		28810	=>	44905,
		28811	=>	44903,
		28812	=>	44900,
		28813	=>	44897,
		28814	=>	44894,
		28815	=>	44891,
		28816	=>	44888,
		28817	=>	44885,
		28818	=>	44882,
		28819	=>	44879,
		28820	=>	44876,
		28821	=>	44873,
		28822	=>	44870,
		28823	=>	44868,
		28824	=>	44865,
		28825	=>	44862,
		28826	=>	44859,
		28827	=>	44856,
		28828	=>	44853,
		28829	=>	44850,
		28830	=>	44847,
		28831	=>	44844,
		28832	=>	44841,
		28833	=>	44838,
		28834	=>	44835,
		28835	=>	44832,
		28836	=>	44830,
		28837	=>	44827,
		28838	=>	44824,
		28839	=>	44821,
		28840	=>	44818,
		28841	=>	44815,
		28842	=>	44812,
		28843	=>	44809,
		28844	=>	44806,
		28845	=>	44803,
		28846	=>	44800,
		28847	=>	44797,
		28848	=>	44794,
		28849	=>	44792,
		28850	=>	44789,
		28851	=>	44786,
		28852	=>	44783,
		28853	=>	44780,
		28854	=>	44777,
		28855	=>	44774,
		28856	=>	44771,
		28857	=>	44768,
		28858	=>	44765,
		28859	=>	44762,
		28860	=>	44759,
		28861	=>	44756,
		28862	=>	44754,
		28863	=>	44751,
		28864	=>	44748,
		28865	=>	44745,
		28866	=>	44742,
		28867	=>	44739,
		28868	=>	44736,
		28869	=>	44733,
		28870	=>	44730,
		28871	=>	44727,
		28872	=>	44724,
		28873	=>	44721,
		28874	=>	44718,
		28875	=>	44716,
		28876	=>	44713,
		28877	=>	44710,
		28878	=>	44707,
		28879	=>	44704,
		28880	=>	44701,
		28881	=>	44698,
		28882	=>	44695,
		28883	=>	44692,
		28884	=>	44689,
		28885	=>	44686,
		28886	=>	44683,
		28887	=>	44680,
		28888	=>	44678,
		28889	=>	44675,
		28890	=>	44672,
		28891	=>	44669,
		28892	=>	44666,
		28893	=>	44663,
		28894	=>	44660,
		28895	=>	44657,
		28896	=>	44654,
		28897	=>	44651,
		28898	=>	44648,
		28899	=>	44645,
		28900	=>	44642,
		28901	=>	44639,
		28902	=>	44637,
		28903	=>	44634,
		28904	=>	44631,
		28905	=>	44628,
		28906	=>	44625,
		28907	=>	44622,
		28908	=>	44619,
		28909	=>	44616,
		28910	=>	44613,
		28911	=>	44610,
		28912	=>	44607,
		28913	=>	44604,
		28914	=>	44601,
		28915	=>	44598,
		28916	=>	44596,
		28917	=>	44593,
		28918	=>	44590,
		28919	=>	44587,
		28920	=>	44584,
		28921	=>	44581,
		28922	=>	44578,
		28923	=>	44575,
		28924	=>	44572,
		28925	=>	44569,
		28926	=>	44566,
		28927	=>	44563,
		28928	=>	44560,
		28929	=>	44557,
		28930	=>	44554,
		28931	=>	44552,
		28932	=>	44549,
		28933	=>	44546,
		28934	=>	44543,
		28935	=>	44540,
		28936	=>	44537,
		28937	=>	44534,
		28938	=>	44531,
		28939	=>	44528,
		28940	=>	44525,
		28941	=>	44522,
		28942	=>	44519,
		28943	=>	44516,
		28944	=>	44513,
		28945	=>	44511,
		28946	=>	44508,
		28947	=>	44505,
		28948	=>	44502,
		28949	=>	44499,
		28950	=>	44496,
		28951	=>	44493,
		28952	=>	44490,
		28953	=>	44487,
		28954	=>	44484,
		28955	=>	44481,
		28956	=>	44478,
		28957	=>	44475,
		28958	=>	44472,
		28959	=>	44469,
		28960	=>	44467,
		28961	=>	44464,
		28962	=>	44461,
		28963	=>	44458,
		28964	=>	44455,
		28965	=>	44452,
		28966	=>	44449,
		28967	=>	44446,
		28968	=>	44443,
		28969	=>	44440,
		28970	=>	44437,
		28971	=>	44434,
		28972	=>	44431,
		28973	=>	44428,
		28974	=>	44425,
		28975	=>	44422,
		28976	=>	44420,
		28977	=>	44417,
		28978	=>	44414,
		28979	=>	44411,
		28980	=>	44408,
		28981	=>	44405,
		28982	=>	44402,
		28983	=>	44399,
		28984	=>	44396,
		28985	=>	44393,
		28986	=>	44390,
		28987	=>	44387,
		28988	=>	44384,
		28989	=>	44381,
		28990	=>	44378,
		28991	=>	44375,
		28992	=>	44373,
		28993	=>	44370,
		28994	=>	44367,
		28995	=>	44364,
		28996	=>	44361,
		28997	=>	44358,
		28998	=>	44355,
		28999	=>	44352,
		29000	=>	44349,
		29001	=>	44346,
		29002	=>	44343,
		29003	=>	44340,
		29004	=>	44337,
		29005	=>	44334,
		29006	=>	44331,
		29007	=>	44328,
		29008	=>	44326,
		29009	=>	44323,
		29010	=>	44320,
		29011	=>	44317,
		29012	=>	44314,
		29013	=>	44311,
		29014	=>	44308,
		29015	=>	44305,
		29016	=>	44302,
		29017	=>	44299,
		29018	=>	44296,
		29019	=>	44293,
		29020	=>	44290,
		29021	=>	44287,
		29022	=>	44284,
		29023	=>	44281,
		29024	=>	44278,
		29025	=>	44276,
		29026	=>	44273,
		29027	=>	44270,
		29028	=>	44267,
		29029	=>	44264,
		29030	=>	44261,
		29031	=>	44258,
		29032	=>	44255,
		29033	=>	44252,
		29034	=>	44249,
		29035	=>	44246,
		29036	=>	44243,
		29037	=>	44240,
		29038	=>	44237,
		29039	=>	44234,
		29040	=>	44231,
		29041	=>	44228,
		29042	=>	44226,
		29043	=>	44223,
		29044	=>	44220,
		29045	=>	44217,
		29046	=>	44214,
		29047	=>	44211,
		29048	=>	44208,
		29049	=>	44205,
		29050	=>	44202,
		29051	=>	44199,
		29052	=>	44196,
		29053	=>	44193,
		29054	=>	44190,
		29055	=>	44187,
		29056	=>	44184,
		29057	=>	44181,
		29058	=>	44178,
		29059	=>	44175,
		29060	=>	44173,
		29061	=>	44170,
		29062	=>	44167,
		29063	=>	44164,
		29064	=>	44161,
		29065	=>	44158,
		29066	=>	44155,
		29067	=>	44152,
		29068	=>	44149,
		29069	=>	44146,
		29070	=>	44143,
		29071	=>	44140,
		29072	=>	44137,
		29073	=>	44134,
		29074	=>	44131,
		29075	=>	44128,
		29076	=>	44125,
		29077	=>	44122,
		29078	=>	44120,
		29079	=>	44117,
		29080	=>	44114,
		29081	=>	44111,
		29082	=>	44108,
		29083	=>	44105,
		29084	=>	44102,
		29085	=>	44099,
		29086	=>	44096,
		29087	=>	44093,
		29088	=>	44090,
		29089	=>	44087,
		29090	=>	44084,
		29091	=>	44081,
		29092	=>	44078,
		29093	=>	44075,
		29094	=>	44072,
		29095	=>	44069,
		29096	=>	44066,
		29097	=>	44063,
		29098	=>	44061,
		29099	=>	44058,
		29100	=>	44055,
		29101	=>	44052,
		29102	=>	44049,
		29103	=>	44046,
		29104	=>	44043,
		29105	=>	44040,
		29106	=>	44037,
		29107	=>	44034,
		29108	=>	44031,
		29109	=>	44028,
		29110	=>	44025,
		29111	=>	44022,
		29112	=>	44019,
		29113	=>	44016,
		29114	=>	44013,
		29115	=>	44010,
		29116	=>	44007,
		29117	=>	44004,
		29118	=>	44002,
		29119	=>	43999,
		29120	=>	43996,
		29121	=>	43993,
		29122	=>	43990,
		29123	=>	43987,
		29124	=>	43984,
		29125	=>	43981,
		29126	=>	43978,
		29127	=>	43975,
		29128	=>	43972,
		29129	=>	43969,
		29130	=>	43966,
		29131	=>	43963,
		29132	=>	43960,
		29133	=>	43957,
		29134	=>	43954,
		29135	=>	43951,
		29136	=>	43948,
		29137	=>	43945,
		29138	=>	43942,
		29139	=>	43940,
		29140	=>	43937,
		29141	=>	43934,
		29142	=>	43931,
		29143	=>	43928,
		29144	=>	43925,
		29145	=>	43922,
		29146	=>	43919,
		29147	=>	43916,
		29148	=>	43913,
		29149	=>	43910,
		29150	=>	43907,
		29151	=>	43904,
		29152	=>	43901,
		29153	=>	43898,
		29154	=>	43895,
		29155	=>	43892,
		29156	=>	43889,
		29157	=>	43886,
		29158	=>	43883,
		29159	=>	43880,
		29160	=>	43877,
		29161	=>	43875,
		29162	=>	43872,
		29163	=>	43869,
		29164	=>	43866,
		29165	=>	43863,
		29166	=>	43860,
		29167	=>	43857,
		29168	=>	43854,
		29169	=>	43851,
		29170	=>	43848,
		29171	=>	43845,
		29172	=>	43842,
		29173	=>	43839,
		29174	=>	43836,
		29175	=>	43833,
		29176	=>	43830,
		29177	=>	43827,
		29178	=>	43824,
		29179	=>	43821,
		29180	=>	43818,
		29181	=>	43815,
		29182	=>	43812,
		29183	=>	43809,
		29184	=>	43807,
		29185	=>	43804,
		29186	=>	43801,
		29187	=>	43798,
		29188	=>	43795,
		29189	=>	43792,
		29190	=>	43789,
		29191	=>	43786,
		29192	=>	43783,
		29193	=>	43780,
		29194	=>	43777,
		29195	=>	43774,
		29196	=>	43771,
		29197	=>	43768,
		29198	=>	43765,
		29199	=>	43762,
		29200	=>	43759,
		29201	=>	43756,
		29202	=>	43753,
		29203	=>	43750,
		29204	=>	43747,
		29205	=>	43744,
		29206	=>	43741,
		29207	=>	43738,
		29208	=>	43736,
		29209	=>	43733,
		29210	=>	43730,
		29211	=>	43727,
		29212	=>	43724,
		29213	=>	43721,
		29214	=>	43718,
		29215	=>	43715,
		29216	=>	43712,
		29217	=>	43709,
		29218	=>	43706,
		29219	=>	43703,
		29220	=>	43700,
		29221	=>	43697,
		29222	=>	43694,
		29223	=>	43691,
		29224	=>	43688,
		29225	=>	43685,
		29226	=>	43682,
		29227	=>	43679,
		29228	=>	43676,
		29229	=>	43673,
		29230	=>	43670,
		29231	=>	43667,
		29232	=>	43664,
		29233	=>	43661,
		29234	=>	43659,
		29235	=>	43656,
		29236	=>	43653,
		29237	=>	43650,
		29238	=>	43647,
		29239	=>	43644,
		29240	=>	43641,
		29241	=>	43638,
		29242	=>	43635,
		29243	=>	43632,
		29244	=>	43629,
		29245	=>	43626,
		29246	=>	43623,
		29247	=>	43620,
		29248	=>	43617,
		29249	=>	43614,
		29250	=>	43611,
		29251	=>	43608,
		29252	=>	43605,
		29253	=>	43602,
		29254	=>	43599,
		29255	=>	43596,
		29256	=>	43593,
		29257	=>	43590,
		29258	=>	43587,
		29259	=>	43584,
		29260	=>	43581,
		29261	=>	43578,
		29262	=>	43576,
		29263	=>	43573,
		29264	=>	43570,
		29265	=>	43567,
		29266	=>	43564,
		29267	=>	43561,
		29268	=>	43558,
		29269	=>	43555,
		29270	=>	43552,
		29271	=>	43549,
		29272	=>	43546,
		29273	=>	43543,
		29274	=>	43540,
		29275	=>	43537,
		29276	=>	43534,
		29277	=>	43531,
		29278	=>	43528,
		29279	=>	43525,
		29280	=>	43522,
		29281	=>	43519,
		29282	=>	43516,
		29283	=>	43513,
		29284	=>	43510,
		29285	=>	43507,
		29286	=>	43504,
		29287	=>	43501,
		29288	=>	43498,
		29289	=>	43495,
		29290	=>	43492,
		29291	=>	43489,
		29292	=>	43486,
		29293	=>	43484,
		29294	=>	43481,
		29295	=>	43478,
		29296	=>	43475,
		29297	=>	43472,
		29298	=>	43469,
		29299	=>	43466,
		29300	=>	43463,
		29301	=>	43460,
		29302	=>	43457,
		29303	=>	43454,
		29304	=>	43451,
		29305	=>	43448,
		29306	=>	43445,
		29307	=>	43442,
		29308	=>	43439,
		29309	=>	43436,
		29310	=>	43433,
		29311	=>	43430,
		29312	=>	43427,
		29313	=>	43424,
		29314	=>	43421,
		29315	=>	43418,
		29316	=>	43415,
		29317	=>	43412,
		29318	=>	43409,
		29319	=>	43406,
		29320	=>	43403,
		29321	=>	43400,
		29322	=>	43397,
		29323	=>	43394,
		29324	=>	43391,
		29325	=>	43388,
		29326	=>	43386,
		29327	=>	43383,
		29328	=>	43380,
		29329	=>	43377,
		29330	=>	43374,
		29331	=>	43371,
		29332	=>	43368,
		29333	=>	43365,
		29334	=>	43362,
		29335	=>	43359,
		29336	=>	43356,
		29337	=>	43353,
		29338	=>	43350,
		29339	=>	43347,
		29340	=>	43344,
		29341	=>	43341,
		29342	=>	43338,
		29343	=>	43335,
		29344	=>	43332,
		29345	=>	43329,
		29346	=>	43326,
		29347	=>	43323,
		29348	=>	43320,
		29349	=>	43317,
		29350	=>	43314,
		29351	=>	43311,
		29352	=>	43308,
		29353	=>	43305,
		29354	=>	43302,
		29355	=>	43299,
		29356	=>	43296,
		29357	=>	43293,
		29358	=>	43290,
		29359	=>	43287,
		29360	=>	43284,
		29361	=>	43281,
		29362	=>	43278,
		29363	=>	43275,
		29364	=>	43272,
		29365	=>	43270,
		29366	=>	43267,
		29367	=>	43264,
		29368	=>	43261,
		29369	=>	43258,
		29370	=>	43255,
		29371	=>	43252,
		29372	=>	43249,
		29373	=>	43246,
		29374	=>	43243,
		29375	=>	43240,
		29376	=>	43237,
		29377	=>	43234,
		29378	=>	43231,
		29379	=>	43228,
		29380	=>	43225,
		29381	=>	43222,
		29382	=>	43219,
		29383	=>	43216,
		29384	=>	43213,
		29385	=>	43210,
		29386	=>	43207,
		29387	=>	43204,
		29388	=>	43201,
		29389	=>	43198,
		29390	=>	43195,
		29391	=>	43192,
		29392	=>	43189,
		29393	=>	43186,
		29394	=>	43183,
		29395	=>	43180,
		29396	=>	43177,
		29397	=>	43174,
		29398	=>	43171,
		29399	=>	43168,
		29400	=>	43165,
		29401	=>	43162,
		29402	=>	43159,
		29403	=>	43156,
		29404	=>	43153,
		29405	=>	43150,
		29406	=>	43147,
		29407	=>	43144,
		29408	=>	43141,
		29409	=>	43138,
		29410	=>	43136,
		29411	=>	43133,
		29412	=>	43130,
		29413	=>	43127,
		29414	=>	43124,
		29415	=>	43121,
		29416	=>	43118,
		29417	=>	43115,
		29418	=>	43112,
		29419	=>	43109,
		29420	=>	43106,
		29421	=>	43103,
		29422	=>	43100,
		29423	=>	43097,
		29424	=>	43094,
		29425	=>	43091,
		29426	=>	43088,
		29427	=>	43085,
		29428	=>	43082,
		29429	=>	43079,
		29430	=>	43076,
		29431	=>	43073,
		29432	=>	43070,
		29433	=>	43067,
		29434	=>	43064,
		29435	=>	43061,
		29436	=>	43058,
		29437	=>	43055,
		29438	=>	43052,
		29439	=>	43049,
		29440	=>	43046,
		29441	=>	43043,
		29442	=>	43040,
		29443	=>	43037,
		29444	=>	43034,
		29445	=>	43031,
		29446	=>	43028,
		29447	=>	43025,
		29448	=>	43022,
		29449	=>	43019,
		29450	=>	43016,
		29451	=>	43013,
		29452	=>	43010,
		29453	=>	43007,
		29454	=>	43004,
		29455	=>	43001,
		29456	=>	42998,
		29457	=>	42995,
		29458	=>	42992,
		29459	=>	42989,
		29460	=>	42986,
		29461	=>	42983,
		29462	=>	42980,
		29463	=>	42977,
		29464	=>	42974,
		29465	=>	42971,
		29466	=>	42968,
		29467	=>	42965,
		29468	=>	42963,
		29469	=>	42960,
		29470	=>	42957,
		29471	=>	42954,
		29472	=>	42951,
		29473	=>	42948,
		29474	=>	42945,
		29475	=>	42942,
		29476	=>	42939,
		29477	=>	42936,
		29478	=>	42933,
		29479	=>	42930,
		29480	=>	42927,
		29481	=>	42924,
		29482	=>	42921,
		29483	=>	42918,
		29484	=>	42915,
		29485	=>	42912,
		29486	=>	42909,
		29487	=>	42906,
		29488	=>	42903,
		29489	=>	42900,
		29490	=>	42897,
		29491	=>	42894,
		29492	=>	42891,
		29493	=>	42888,
		29494	=>	42885,
		29495	=>	42882,
		29496	=>	42879,
		29497	=>	42876,
		29498	=>	42873,
		29499	=>	42870,
		29500	=>	42867,
		29501	=>	42864,
		29502	=>	42861,
		29503	=>	42858,
		29504	=>	42855,
		29505	=>	42852,
		29506	=>	42849,
		29507	=>	42846,
		29508	=>	42843,
		29509	=>	42840,
		29510	=>	42837,
		29511	=>	42834,
		29512	=>	42831,
		29513	=>	42828,
		29514	=>	42825,
		29515	=>	42822,
		29516	=>	42819,
		29517	=>	42816,
		29518	=>	42813,
		29519	=>	42810,
		29520	=>	42807,
		29521	=>	42804,
		29522	=>	42801,
		29523	=>	42798,
		29524	=>	42795,
		29525	=>	42792,
		29526	=>	42789,
		29527	=>	42786,
		29528	=>	42783,
		29529	=>	42780,
		29530	=>	42777,
		29531	=>	42774,
		29532	=>	42771,
		29533	=>	42768,
		29534	=>	42765,
		29535	=>	42762,
		29536	=>	42759,
		29537	=>	42756,
		29538	=>	42753,
		29539	=>	42750,
		29540	=>	42747,
		29541	=>	42744,
		29542	=>	42741,
		29543	=>	42738,
		29544	=>	42735,
		29545	=>	42732,
		29546	=>	42729,
		29547	=>	42726,
		29548	=>	42723,
		29549	=>	42720,
		29550	=>	42717,
		29551	=>	42714,
		29552	=>	42711,
		29553	=>	42708,
		29554	=>	42705,
		29555	=>	42702,
		29556	=>	42699,
		29557	=>	42696,
		29558	=>	42693,
		29559	=>	42690,
		29560	=>	42687,
		29561	=>	42684,
		29562	=>	42681,
		29563	=>	42678,
		29564	=>	42675,
		29565	=>	42672,
		29566	=>	42669,
		29567	=>	42666,
		29568	=>	42663,
		29569	=>	42660,
		29570	=>	42657,
		29571	=>	42654,
		29572	=>	42651,
		29573	=>	42649,
		29574	=>	42646,
		29575	=>	42643,
		29576	=>	42640,
		29577	=>	42637,
		29578	=>	42634,
		29579	=>	42631,
		29580	=>	42628,
		29581	=>	42625,
		29582	=>	42622,
		29583	=>	42619,
		29584	=>	42616,
		29585	=>	42613,
		29586	=>	42610,
		29587	=>	42607,
		29588	=>	42604,
		29589	=>	42601,
		29590	=>	42598,
		29591	=>	42595,
		29592	=>	42592,
		29593	=>	42589,
		29594	=>	42586,
		29595	=>	42583,
		29596	=>	42580,
		29597	=>	42577,
		29598	=>	42574,
		29599	=>	42571,
		29600	=>	42568,
		29601	=>	42565,
		29602	=>	42562,
		29603	=>	42559,
		29604	=>	42556,
		29605	=>	42553,
		29606	=>	42550,
		29607	=>	42547,
		29608	=>	42544,
		29609	=>	42541,
		29610	=>	42538,
		29611	=>	42535,
		29612	=>	42532,
		29613	=>	42529,
		29614	=>	42526,
		29615	=>	42523,
		29616	=>	42520,
		29617	=>	42517,
		29618	=>	42514,
		29619	=>	42511,
		29620	=>	42508,
		29621	=>	42505,
		29622	=>	42502,
		29623	=>	42499,
		29624	=>	42496,
		29625	=>	42493,
		29626	=>	42490,
		29627	=>	42487,
		29628	=>	42484,
		29629	=>	42481,
		29630	=>	42478,
		29631	=>	42475,
		29632	=>	42472,
		29633	=>	42469,
		29634	=>	42466,
		29635	=>	42463,
		29636	=>	42460,
		29637	=>	42457,
		29638	=>	42454,
		29639	=>	42451,
		29640	=>	42448,
		29641	=>	42445,
		29642	=>	42442,
		29643	=>	42439,
		29644	=>	42436,
		29645	=>	42433,
		29646	=>	42430,
		29647	=>	42427,
		29648	=>	42424,
		29649	=>	42421,
		29650	=>	42418,
		29651	=>	42415,
		29652	=>	42412,
		29653	=>	42409,
		29654	=>	42406,
		29655	=>	42403,
		29656	=>	42400,
		29657	=>	42397,
		29658	=>	42394,
		29659	=>	42391,
		29660	=>	42388,
		29661	=>	42385,
		29662	=>	42382,
		29663	=>	42379,
		29664	=>	42376,
		29665	=>	42373,
		29666	=>	42370,
		29667	=>	42367,
		29668	=>	42364,
		29669	=>	42361,
		29670	=>	42358,
		29671	=>	42355,
		29672	=>	42352,
		29673	=>	42349,
		29674	=>	42346,
		29675	=>	42343,
		29676	=>	42340,
		29677	=>	42337,
		29678	=>	42334,
		29679	=>	42330,
		29680	=>	42327,
		29681	=>	42324,
		29682	=>	42321,
		29683	=>	42318,
		29684	=>	42315,
		29685	=>	42312,
		29686	=>	42309,
		29687	=>	42306,
		29688	=>	42303,
		29689	=>	42300,
		29690	=>	42297,
		29691	=>	42294,
		29692	=>	42291,
		29693	=>	42288,
		29694	=>	42285,
		29695	=>	42282,
		29696	=>	42279,
		29697	=>	42276,
		29698	=>	42273,
		29699	=>	42270,
		29700	=>	42267,
		29701	=>	42264,
		29702	=>	42261,
		29703	=>	42258,
		29704	=>	42255,
		29705	=>	42252,
		29706	=>	42249,
		29707	=>	42246,
		29708	=>	42243,
		29709	=>	42240,
		29710	=>	42237,
		29711	=>	42234,
		29712	=>	42231,
		29713	=>	42228,
		29714	=>	42225,
		29715	=>	42222,
		29716	=>	42219,
		29717	=>	42216,
		29718	=>	42213,
		29719	=>	42210,
		29720	=>	42207,
		29721	=>	42204,
		29722	=>	42201,
		29723	=>	42198,
		29724	=>	42195,
		29725	=>	42192,
		29726	=>	42189,
		29727	=>	42186,
		29728	=>	42183,
		29729	=>	42180,
		29730	=>	42177,
		29731	=>	42174,
		29732	=>	42171,
		29733	=>	42168,
		29734	=>	42165,
		29735	=>	42162,
		29736	=>	42159,
		29737	=>	42156,
		29738	=>	42153,
		29739	=>	42150,
		29740	=>	42147,
		29741	=>	42144,
		29742	=>	42141,
		29743	=>	42138,
		29744	=>	42135,
		29745	=>	42132,
		29746	=>	42129,
		29747	=>	42126,
		29748	=>	42123,
		29749	=>	42120,
		29750	=>	42117,
		29751	=>	42114,
		29752	=>	42111,
		29753	=>	42108,
		29754	=>	42105,
		29755	=>	42102,
		29756	=>	42099,
		29757	=>	42096,
		29758	=>	42093,
		29759	=>	42090,
		29760	=>	42087,
		29761	=>	42084,
		29762	=>	42081,
		29763	=>	42078,
		29764	=>	42075,
		29765	=>	42072,
		29766	=>	42069,
		29767	=>	42066,
		29768	=>	42063,
		29769	=>	42060,
		29770	=>	42057,
		29771	=>	42054,
		29772	=>	42051,
		29773	=>	42048,
		29774	=>	42045,
		29775	=>	42042,
		29776	=>	42039,
		29777	=>	42036,
		29778	=>	42033,
		29779	=>	42030,
		29780	=>	42027,
		29781	=>	42024,
		29782	=>	42021,
		29783	=>	42018,
		29784	=>	42015,
		29785	=>	42012,
		29786	=>	42008,
		29787	=>	42005,
		29788	=>	42002,
		29789	=>	41999,
		29790	=>	41996,
		29791	=>	41993,
		29792	=>	41990,
		29793	=>	41987,
		29794	=>	41984,
		29795	=>	41981,
		29796	=>	41978,
		29797	=>	41975,
		29798	=>	41972,
		29799	=>	41969,
		29800	=>	41966,
		29801	=>	41963,
		29802	=>	41960,
		29803	=>	41957,
		29804	=>	41954,
		29805	=>	41951,
		29806	=>	41948,
		29807	=>	41945,
		29808	=>	41942,
		29809	=>	41939,
		29810	=>	41936,
		29811	=>	41933,
		29812	=>	41930,
		29813	=>	41927,
		29814	=>	41924,
		29815	=>	41921,
		29816	=>	41918,
		29817	=>	41915,
		29818	=>	41912,
		29819	=>	41909,
		29820	=>	41906,
		29821	=>	41903,
		29822	=>	41900,
		29823	=>	41897,
		29824	=>	41894,
		29825	=>	41891,
		29826	=>	41888,
		29827	=>	41885,
		29828	=>	41882,
		29829	=>	41879,
		29830	=>	41876,
		29831	=>	41873,
		29832	=>	41870,
		29833	=>	41867,
		29834	=>	41864,
		29835	=>	41861,
		29836	=>	41858,
		29837	=>	41855,
		29838	=>	41852,
		29839	=>	41849,
		29840	=>	41846,
		29841	=>	41843,
		29842	=>	41840,
		29843	=>	41837,
		29844	=>	41834,
		29845	=>	41831,
		29846	=>	41827,
		29847	=>	41824,
		29848	=>	41821,
		29849	=>	41818,
		29850	=>	41815,
		29851	=>	41812,
		29852	=>	41809,
		29853	=>	41806,
		29854	=>	41803,
		29855	=>	41800,
		29856	=>	41797,
		29857	=>	41794,
		29858	=>	41791,
		29859	=>	41788,
		29860	=>	41785,
		29861	=>	41782,
		29862	=>	41779,
		29863	=>	41776,
		29864	=>	41773,
		29865	=>	41770,
		29866	=>	41767,
		29867	=>	41764,
		29868	=>	41761,
		29869	=>	41758,
		29870	=>	41755,
		29871	=>	41752,
		29872	=>	41749,
		29873	=>	41746,
		29874	=>	41743,
		29875	=>	41740,
		29876	=>	41737,
		29877	=>	41734,
		29878	=>	41731,
		29879	=>	41728,
		29880	=>	41725,
		29881	=>	41722,
		29882	=>	41719,
		29883	=>	41716,
		29884	=>	41713,
		29885	=>	41710,
		29886	=>	41707,
		29887	=>	41704,
		29888	=>	41701,
		29889	=>	41698,
		29890	=>	41695,
		29891	=>	41692,
		29892	=>	41689,
		29893	=>	41686,
		29894	=>	41682,
		29895	=>	41679,
		29896	=>	41676,
		29897	=>	41673,
		29898	=>	41670,
		29899	=>	41667,
		29900	=>	41664,
		29901	=>	41661,
		29902	=>	41658,
		29903	=>	41655,
		29904	=>	41652,
		29905	=>	41649,
		29906	=>	41646,
		29907	=>	41643,
		29908	=>	41640,
		29909	=>	41637,
		29910	=>	41634,
		29911	=>	41631,
		29912	=>	41628,
		29913	=>	41625,
		29914	=>	41622,
		29915	=>	41619,
		29916	=>	41616,
		29917	=>	41613,
		29918	=>	41610,
		29919	=>	41607,
		29920	=>	41604,
		29921	=>	41601,
		29922	=>	41598,
		29923	=>	41595,
		29924	=>	41592,
		29925	=>	41589,
		29926	=>	41586,
		29927	=>	41583,
		29928	=>	41580,
		29929	=>	41577,
		29930	=>	41574,
		29931	=>	41571,
		29932	=>	41568,
		29933	=>	41565,
		29934	=>	41561,
		29935	=>	41558,
		29936	=>	41555,
		29937	=>	41552,
		29938	=>	41549,
		29939	=>	41546,
		29940	=>	41543,
		29941	=>	41540,
		29942	=>	41537,
		29943	=>	41534,
		29944	=>	41531,
		29945	=>	41528,
		29946	=>	41525,
		29947	=>	41522,
		29948	=>	41519,
		29949	=>	41516,
		29950	=>	41513,
		29951	=>	41510,
		29952	=>	41507,
		29953	=>	41504,
		29954	=>	41501,
		29955	=>	41498,
		29956	=>	41495,
		29957	=>	41492,
		29958	=>	41489,
		29959	=>	41486,
		29960	=>	41483,
		29961	=>	41480,
		29962	=>	41477,
		29963	=>	41474,
		29964	=>	41471,
		29965	=>	41468,
		29966	=>	41465,
		29967	=>	41462,
		29968	=>	41459,
		29969	=>	41456,
		29970	=>	41452,
		29971	=>	41449,
		29972	=>	41446,
		29973	=>	41443,
		29974	=>	41440,
		29975	=>	41437,
		29976	=>	41434,
		29977	=>	41431,
		29978	=>	41428,
		29979	=>	41425,
		29980	=>	41422,
		29981	=>	41419,
		29982	=>	41416,
		29983	=>	41413,
		29984	=>	41410,
		29985	=>	41407,
		29986	=>	41404,
		29987	=>	41401,
		29988	=>	41398,
		29989	=>	41395,
		29990	=>	41392,
		29991	=>	41389,
		29992	=>	41386,
		29993	=>	41383,
		29994	=>	41380,
		29995	=>	41377,
		29996	=>	41374,
		29997	=>	41371,
		29998	=>	41368,
		29999	=>	41365,
		30000	=>	41362,
		30001	=>	41359,
		30002	=>	41356,
		30003	=>	41352,
		30004	=>	41349,
		30005	=>	41346,
		30006	=>	41343,
		30007	=>	41340,
		30008	=>	41337,
		30009	=>	41334,
		30010	=>	41331,
		30011	=>	41328,
		30012	=>	41325,
		30013	=>	41322,
		30014	=>	41319,
		30015	=>	41316,
		30016	=>	41313,
		30017	=>	41310,
		30018	=>	41307,
		30019	=>	41304,
		30020	=>	41301,
		30021	=>	41298,
		30022	=>	41295,
		30023	=>	41292,
		30024	=>	41289,
		30025	=>	41286,
		30026	=>	41283,
		30027	=>	41280,
		30028	=>	41277,
		30029	=>	41274,
		30030	=>	41271,
		30031	=>	41268,
		30032	=>	41265,
		30033	=>	41262,
		30034	=>	41258,
		30035	=>	41255,
		30036	=>	41252,
		30037	=>	41249,
		30038	=>	41246,
		30039	=>	41243,
		30040	=>	41240,
		30041	=>	41237,
		30042	=>	41234,
		30043	=>	41231,
		30044	=>	41228,
		30045	=>	41225,
		30046	=>	41222,
		30047	=>	41219,
		30048	=>	41216,
		30049	=>	41213,
		30050	=>	41210,
		30051	=>	41207,
		30052	=>	41204,
		30053	=>	41201,
		30054	=>	41198,
		30055	=>	41195,
		30056	=>	41192,
		30057	=>	41189,
		30058	=>	41186,
		30059	=>	41183,
		30060	=>	41180,
		30061	=>	41177,
		30062	=>	41173,
		30063	=>	41170,
		30064	=>	41167,
		30065	=>	41164,
		30066	=>	41161,
		30067	=>	41158,
		30068	=>	41155,
		30069	=>	41152,
		30070	=>	41149,
		30071	=>	41146,
		30072	=>	41143,
		30073	=>	41140,
		30074	=>	41137,
		30075	=>	41134,
		30076	=>	41131,
		30077	=>	41128,
		30078	=>	41125,
		30079	=>	41122,
		30080	=>	41119,
		30081	=>	41116,
		30082	=>	41113,
		30083	=>	41110,
		30084	=>	41107,
		30085	=>	41104,
		30086	=>	41101,
		30087	=>	41098,
		30088	=>	41095,
		30089	=>	41091,
		30090	=>	41088,
		30091	=>	41085,
		30092	=>	41082,
		30093	=>	41079,
		30094	=>	41076,
		30095	=>	41073,
		30096	=>	41070,
		30097	=>	41067,
		30098	=>	41064,
		30099	=>	41061,
		30100	=>	41058,
		30101	=>	41055,
		30102	=>	41052,
		30103	=>	41049,
		30104	=>	41046,
		30105	=>	41043,
		30106	=>	41040,
		30107	=>	41037,
		30108	=>	41034,
		30109	=>	41031,
		30110	=>	41028,
		30111	=>	41025,
		30112	=>	41022,
		30113	=>	41019,
		30114	=>	41015,
		30115	=>	41012,
		30116	=>	41009,
		30117	=>	41006,
		30118	=>	41003,
		30119	=>	41000,
		30120	=>	40997,
		30121	=>	40994,
		30122	=>	40991,
		30123	=>	40988,
		30124	=>	40985,
		30125	=>	40982,
		30126	=>	40979,
		30127	=>	40976,
		30128	=>	40973,
		30129	=>	40970,
		30130	=>	40967,
		30131	=>	40964,
		30132	=>	40961,
		30133	=>	40958,
		30134	=>	40955,
		30135	=>	40952,
		30136	=>	40949,
		30137	=>	40946,
		30138	=>	40942,
		30139	=>	40939,
		30140	=>	40936,
		30141	=>	40933,
		30142	=>	40930,
		30143	=>	40927,
		30144	=>	40924,
		30145	=>	40921,
		30146	=>	40918,
		30147	=>	40915,
		30148	=>	40912,
		30149	=>	40909,
		30150	=>	40906,
		30151	=>	40903,
		30152	=>	40900,
		30153	=>	40897,
		30154	=>	40894,
		30155	=>	40891,
		30156	=>	40888,
		30157	=>	40885,
		30158	=>	40882,
		30159	=>	40879,
		30160	=>	40876,
		30161	=>	40872,
		30162	=>	40869,
		30163	=>	40866,
		30164	=>	40863,
		30165	=>	40860,
		30166	=>	40857,
		30167	=>	40854,
		30168	=>	40851,
		30169	=>	40848,
		30170	=>	40845,
		30171	=>	40842,
		30172	=>	40839,
		30173	=>	40836,
		30174	=>	40833,
		30175	=>	40830,
		30176	=>	40827,
		30177	=>	40824,
		30178	=>	40821,
		30179	=>	40818,
		30180	=>	40815,
		30181	=>	40812,
		30182	=>	40809,
		30183	=>	40806,
		30184	=>	40802,
		30185	=>	40799,
		30186	=>	40796,
		30187	=>	40793,
		30188	=>	40790,
		30189	=>	40787,
		30190	=>	40784,
		30191	=>	40781,
		30192	=>	40778,
		30193	=>	40775,
		30194	=>	40772,
		30195	=>	40769,
		30196	=>	40766,
		30197	=>	40763,
		30198	=>	40760,
		30199	=>	40757,
		30200	=>	40754,
		30201	=>	40751,
		30202	=>	40748,
		30203	=>	40745,
		30204	=>	40742,
		30205	=>	40738,
		30206	=>	40735,
		30207	=>	40732,
		30208	=>	40729,
		30209	=>	40726,
		30210	=>	40723,
		30211	=>	40720,
		30212	=>	40717,
		30213	=>	40714,
		30214	=>	40711,
		30215	=>	40708,
		30216	=>	40705,
		30217	=>	40702,
		30218	=>	40699,
		30219	=>	40696,
		30220	=>	40693,
		30221	=>	40690,
		30222	=>	40687,
		30223	=>	40684,
		30224	=>	40681,
		30225	=>	40678,
		30226	=>	40674,
		30227	=>	40671,
		30228	=>	40668,
		30229	=>	40665,
		30230	=>	40662,
		30231	=>	40659,
		30232	=>	40656,
		30233	=>	40653,
		30234	=>	40650,
		30235	=>	40647,
		30236	=>	40644,
		30237	=>	40641,
		30238	=>	40638,
		30239	=>	40635,
		30240	=>	40632,
		30241	=>	40629,
		30242	=>	40626,
		30243	=>	40623,
		30244	=>	40620,
		30245	=>	40617,
		30246	=>	40613,
		30247	=>	40610,
		30248	=>	40607,
		30249	=>	40604,
		30250	=>	40601,
		30251	=>	40598,
		30252	=>	40595,
		30253	=>	40592,
		30254	=>	40589,
		30255	=>	40586,
		30256	=>	40583,
		30257	=>	40580,
		30258	=>	40577,
		30259	=>	40574,
		30260	=>	40571,
		30261	=>	40568,
		30262	=>	40565,
		30263	=>	40562,
		30264	=>	40559,
		30265	=>	40556,
		30266	=>	40552,
		30267	=>	40549,
		30268	=>	40546,
		30269	=>	40543,
		30270	=>	40540,
		30271	=>	40537,
		30272	=>	40534,
		30273	=>	40531,
		30274	=>	40528,
		30275	=>	40525,
		30276	=>	40522,
		30277	=>	40519,
		30278	=>	40516,
		30279	=>	40513,
		30280	=>	40510,
		30281	=>	40507,
		30282	=>	40504,
		30283	=>	40501,
		30284	=>	40498,
		30285	=>	40494,
		30286	=>	40491,
		30287	=>	40488,
		30288	=>	40485,
		30289	=>	40482,
		30290	=>	40479,
		30291	=>	40476,
		30292	=>	40473,
		30293	=>	40470,
		30294	=>	40467,
		30295	=>	40464,
		30296	=>	40461,
		30297	=>	40458,
		30298	=>	40455,
		30299	=>	40452,
		30300	=>	40449,
		30301	=>	40446,
		30302	=>	40443,
		30303	=>	40440,
		30304	=>	40436,
		30305	=>	40433,
		30306	=>	40430,
		30307	=>	40427,
		30308	=>	40424,
		30309	=>	40421,
		30310	=>	40418,
		30311	=>	40415,
		30312	=>	40412,
		30313	=>	40409,
		30314	=>	40406,
		30315	=>	40403,
		30316	=>	40400,
		30317	=>	40397,
		30318	=>	40394,
		30319	=>	40391,
		30320	=>	40388,
		30321	=>	40385,
		30322	=>	40381,
		30323	=>	40378,
		30324	=>	40375,
		30325	=>	40372,
		30326	=>	40369,
		30327	=>	40366,
		30328	=>	40363,
		30329	=>	40360,
		30330	=>	40357,
		30331	=>	40354,
		30332	=>	40351,
		30333	=>	40348,
		30334	=>	40345,
		30335	=>	40342,
		30336	=>	40339,
		30337	=>	40336,
		30338	=>	40333,
		30339	=>	40330,
		30340	=>	40326,
		30341	=>	40323,
		30342	=>	40320,
		30343	=>	40317,
		30344	=>	40314,
		30345	=>	40311,
		30346	=>	40308,
		30347	=>	40305,
		30348	=>	40302,
		30349	=>	40299,
		30350	=>	40296,
		30351	=>	40293,
		30352	=>	40290,
		30353	=>	40287,
		30354	=>	40284,
		30355	=>	40281,
		30356	=>	40278,
		30357	=>	40274,
		30358	=>	40271,
		30359	=>	40268,
		30360	=>	40265,
		30361	=>	40262,
		30362	=>	40259,
		30363	=>	40256,
		30364	=>	40253,
		30365	=>	40250,
		30366	=>	40247,
		30367	=>	40244,
		30368	=>	40241,
		30369	=>	40238,
		30370	=>	40235,
		30371	=>	40232,
		30372	=>	40229,
		30373	=>	40226,
		30374	=>	40222,
		30375	=>	40219,
		30376	=>	40216,
		30377	=>	40213,
		30378	=>	40210,
		30379	=>	40207,
		30380	=>	40204,
		30381	=>	40201,
		30382	=>	40198,
		30383	=>	40195,
		30384	=>	40192,
		30385	=>	40189,
		30386	=>	40186,
		30387	=>	40183,
		30388	=>	40180,
		30389	=>	40177,
		30390	=>	40174,
		30391	=>	40170,
		30392	=>	40167,
		30393	=>	40164,
		30394	=>	40161,
		30395	=>	40158,
		30396	=>	40155,
		30397	=>	40152,
		30398	=>	40149,
		30399	=>	40146,
		30400	=>	40143,
		30401	=>	40140,
		30402	=>	40137,
		30403	=>	40134,
		30404	=>	40131,
		30405	=>	40128,
		30406	=>	40125,
		30407	=>	40122,
		30408	=>	40118,
		30409	=>	40115,
		30410	=>	40112,
		30411	=>	40109,
		30412	=>	40106,
		30413	=>	40103,
		30414	=>	40100,
		30415	=>	40097,
		30416	=>	40094,
		30417	=>	40091,
		30418	=>	40088,
		30419	=>	40085,
		30420	=>	40082,
		30421	=>	40079,
		30422	=>	40076,
		30423	=>	40073,
		30424	=>	40069,
		30425	=>	40066,
		30426	=>	40063,
		30427	=>	40060,
		30428	=>	40057,
		30429	=>	40054,
		30430	=>	40051,
		30431	=>	40048,
		30432	=>	40045,
		30433	=>	40042,
		30434	=>	40039,
		30435	=>	40036,
		30436	=>	40033,
		30437	=>	40030,
		30438	=>	40027,
		30439	=>	40024,
		30440	=>	40020,
		30441	=>	40017,
		30442	=>	40014,
		30443	=>	40011,
		30444	=>	40008,
		30445	=>	40005,
		30446	=>	40002,
		30447	=>	39999,
		30448	=>	39996,
		30449	=>	39993,
		30450	=>	39990,
		30451	=>	39987,
		30452	=>	39984,
		30453	=>	39981,
		30454	=>	39978,
		30455	=>	39974,
		30456	=>	39971,
		30457	=>	39968,
		30458	=>	39965,
		30459	=>	39962,
		30460	=>	39959,
		30461	=>	39956,
		30462	=>	39953,
		30463	=>	39950,
		30464	=>	39947,
		30465	=>	39944,
		30466	=>	39941,
		30467	=>	39938,
		30468	=>	39935,
		30469	=>	39932,
		30470	=>	39929,
		30471	=>	39925,
		30472	=>	39922,
		30473	=>	39919,
		30474	=>	39916,
		30475	=>	39913,
		30476	=>	39910,
		30477	=>	39907,
		30478	=>	39904,
		30479	=>	39901,
		30480	=>	39898,
		30481	=>	39895,
		30482	=>	39892,
		30483	=>	39889,
		30484	=>	39886,
		30485	=>	39883,
		30486	=>	39879,
		30487	=>	39876,
		30488	=>	39873,
		30489	=>	39870,
		30490	=>	39867,
		30491	=>	39864,
		30492	=>	39861,
		30493	=>	39858,
		30494	=>	39855,
		30495	=>	39852,
		30496	=>	39849,
		30497	=>	39846,
		30498	=>	39843,
		30499	=>	39840,
		30500	=>	39837,
		30501	=>	39833,
		30502	=>	39830,
		30503	=>	39827,
		30504	=>	39824,
		30505	=>	39821,
		30506	=>	39818,
		30507	=>	39815,
		30508	=>	39812,
		30509	=>	39809,
		30510	=>	39806,
		30511	=>	39803,
		30512	=>	39800,
		30513	=>	39797,
		30514	=>	39794,
		30515	=>	39790,
		30516	=>	39787,
		30517	=>	39784,
		30518	=>	39781,
		30519	=>	39778,
		30520	=>	39775,
		30521	=>	39772,
		30522	=>	39769,
		30523	=>	39766,
		30524	=>	39763,
		30525	=>	39760,
		30526	=>	39757,
		30527	=>	39754,
		30528	=>	39751,
		30529	=>	39748,
		30530	=>	39744,
		30531	=>	39741,
		30532	=>	39738,
		30533	=>	39735,
		30534	=>	39732,
		30535	=>	39729,
		30536	=>	39726,
		30537	=>	39723,
		30538	=>	39720,
		30539	=>	39717,
		30540	=>	39714,
		30541	=>	39711,
		30542	=>	39708,
		30543	=>	39705,
		30544	=>	39701,
		30545	=>	39698,
		30546	=>	39695,
		30547	=>	39692,
		30548	=>	39689,
		30549	=>	39686,
		30550	=>	39683,
		30551	=>	39680,
		30552	=>	39677,
		30553	=>	39674,
		30554	=>	39671,
		30555	=>	39668,
		30556	=>	39665,
		30557	=>	39662,
		30558	=>	39658,
		30559	=>	39655,
		30560	=>	39652,
		30561	=>	39649,
		30562	=>	39646,
		30563	=>	39643,
		30564	=>	39640,
		30565	=>	39637,
		30566	=>	39634,
		30567	=>	39631,
		30568	=>	39628,
		30569	=>	39625,
		30570	=>	39622,
		30571	=>	39619,
		30572	=>	39615,
		30573	=>	39612,
		30574	=>	39609,
		30575	=>	39606,
		30576	=>	39603,
		30577	=>	39600,
		30578	=>	39597,
		30579	=>	39594,
		30580	=>	39591,
		30581	=>	39588,
		30582	=>	39585,
		30583	=>	39582,
		30584	=>	39579,
		30585	=>	39576,
		30586	=>	39572,
		30587	=>	39569,
		30588	=>	39566,
		30589	=>	39563,
		30590	=>	39560,
		30591	=>	39557,
		30592	=>	39554,
		30593	=>	39551,
		30594	=>	39548,
		30595	=>	39545,
		30596	=>	39542,
		30597	=>	39539,
		30598	=>	39536,
		30599	=>	39533,
		30600	=>	39529,
		30601	=>	39526,
		30602	=>	39523,
		30603	=>	39520,
		30604	=>	39517,
		30605	=>	39514,
		30606	=>	39511,
		30607	=>	39508,
		30608	=>	39505,
		30609	=>	39502,
		30610	=>	39499,
		30611	=>	39496,
		30612	=>	39493,
		30613	=>	39489,
		30614	=>	39486,
		30615	=>	39483,
		30616	=>	39480,
		30617	=>	39477,
		30618	=>	39474,
		30619	=>	39471,
		30620	=>	39468,
		30621	=>	39465,
		30622	=>	39462,
		30623	=>	39459,
		30624	=>	39456,
		30625	=>	39453,
		30626	=>	39449,
		30627	=>	39446,
		30628	=>	39443,
		30629	=>	39440,
		30630	=>	39437,
		30631	=>	39434,
		30632	=>	39431,
		30633	=>	39428,
		30634	=>	39425,
		30635	=>	39422,
		30636	=>	39419,
		30637	=>	39416,
		30638	=>	39413,
		30639	=>	39410,
		30640	=>	39406,
		30641	=>	39403,
		30642	=>	39400,
		30643	=>	39397,
		30644	=>	39394,
		30645	=>	39391,
		30646	=>	39388,
		30647	=>	39385,
		30648	=>	39382,
		30649	=>	39379,
		30650	=>	39376,
		30651	=>	39373,
		30652	=>	39370,
		30653	=>	39366,
		30654	=>	39363,
		30655	=>	39360,
		30656	=>	39357,
		30657	=>	39354,
		30658	=>	39351,
		30659	=>	39348,
		30660	=>	39345,
		30661	=>	39342,
		30662	=>	39339,
		30663	=>	39336,
		30664	=>	39333,
		30665	=>	39329,
		30666	=>	39326,
		30667	=>	39323,
		30668	=>	39320,
		30669	=>	39317,
		30670	=>	39314,
		30671	=>	39311,
		30672	=>	39308,
		30673	=>	39305,
		30674	=>	39302,
		30675	=>	39299,
		30676	=>	39296,
		30677	=>	39293,
		30678	=>	39289,
		30679	=>	39286,
		30680	=>	39283,
		30681	=>	39280,
		30682	=>	39277,
		30683	=>	39274,
		30684	=>	39271,
		30685	=>	39268,
		30686	=>	39265,
		30687	=>	39262,
		30688	=>	39259,
		30689	=>	39256,
		30690	=>	39253,
		30691	=>	39249,
		30692	=>	39246,
		30693	=>	39243,
		30694	=>	39240,
		30695	=>	39237,
		30696	=>	39234,
		30697	=>	39231,
		30698	=>	39228,
		30699	=>	39225,
		30700	=>	39222,
		30701	=>	39219,
		30702	=>	39216,
		30703	=>	39212,
		30704	=>	39209,
		30705	=>	39206,
		30706	=>	39203,
		30707	=>	39200,
		30708	=>	39197,
		30709	=>	39194,
		30710	=>	39191,
		30711	=>	39188,
		30712	=>	39185,
		30713	=>	39182,
		30714	=>	39179,
		30715	=>	39176,
		30716	=>	39172,
		30717	=>	39169,
		30718	=>	39166,
		30719	=>	39163,
		30720	=>	39160,
		30721	=>	39157,
		30722	=>	39154,
		30723	=>	39151,
		30724	=>	39148,
		30725	=>	39145,
		30726	=>	39142,
		30727	=>	39139,
		30728	=>	39135,
		30729	=>	39132,
		30730	=>	39129,
		30731	=>	39126,
		30732	=>	39123,
		30733	=>	39120,
		30734	=>	39117,
		30735	=>	39114,
		30736	=>	39111,
		30737	=>	39108,
		30738	=>	39105,
		30739	=>	39102,
		30740	=>	39098,
		30741	=>	39095,
		30742	=>	39092,
		30743	=>	39089,
		30744	=>	39086,
		30745	=>	39083,
		30746	=>	39080,
		30747	=>	39077,
		30748	=>	39074,
		30749	=>	39071,
		30750	=>	39068,
		30751	=>	39065,
		30752	=>	39061,
		30753	=>	39058,
		30754	=>	39055,
		30755	=>	39052,
		30756	=>	39049,
		30757	=>	39046,
		30758	=>	39043,
		30759	=>	39040,
		30760	=>	39037,
		30761	=>	39034,
		30762	=>	39031,
		30763	=>	39028,
		30764	=>	39024,
		30765	=>	39021,
		30766	=>	39018,
		30767	=>	39015,
		30768	=>	39012,
		30769	=>	39009,
		30770	=>	39006,
		30771	=>	39003,
		30772	=>	39000,
		30773	=>	38997,
		30774	=>	38994,
		30775	=>	38991,
		30776	=>	38987,
		30777	=>	38984,
		30778	=>	38981,
		30779	=>	38978,
		30780	=>	38975,
		30781	=>	38972,
		30782	=>	38969,
		30783	=>	38966,
		30784	=>	38963,
		30785	=>	38960,
		30786	=>	38957,
		30787	=>	38954,
		30788	=>	38950,
		30789	=>	38947,
		30790	=>	38944,
		30791	=>	38941,
		30792	=>	38938,
		30793	=>	38935,
		30794	=>	38932,
		30795	=>	38929,
		30796	=>	38926,
		30797	=>	38923,
		30798	=>	38920,
		30799	=>	38917,
		30800	=>	38913,
		30801	=>	38910,
		30802	=>	38907,
		30803	=>	38904,
		30804	=>	38901,
		30805	=>	38898,
		30806	=>	38895,
		30807	=>	38892,
		30808	=>	38889,
		30809	=>	38886,
		30810	=>	38883,
		30811	=>	38879,
		30812	=>	38876,
		30813	=>	38873,
		30814	=>	38870,
		30815	=>	38867,
		30816	=>	38864,
		30817	=>	38861,
		30818	=>	38858,
		30819	=>	38855,
		30820	=>	38852,
		30821	=>	38849,
		30822	=>	38846,
		30823	=>	38842,
		30824	=>	38839,
		30825	=>	38836,
		30826	=>	38833,
		30827	=>	38830,
		30828	=>	38827,
		30829	=>	38824,
		30830	=>	38821,
		30831	=>	38818,
		30832	=>	38815,
		30833	=>	38812,
		30834	=>	38808,
		30835	=>	38805,
		30836	=>	38802,
		30837	=>	38799,
		30838	=>	38796,
		30839	=>	38793,
		30840	=>	38790,
		30841	=>	38787,
		30842	=>	38784,
		30843	=>	38781,
		30844	=>	38778,
		30845	=>	38775,
		30846	=>	38771,
		30847	=>	38768,
		30848	=>	38765,
		30849	=>	38762,
		30850	=>	38759,
		30851	=>	38756,
		30852	=>	38753,
		30853	=>	38750,
		30854	=>	38747,
		30855	=>	38744,
		30856	=>	38741,
		30857	=>	38737,
		30858	=>	38734,
		30859	=>	38731,
		30860	=>	38728,
		30861	=>	38725,
		30862	=>	38722,
		30863	=>	38719,
		30864	=>	38716,
		30865	=>	38713,
		30866	=>	38710,
		30867	=>	38707,
		30868	=>	38703,
		30869	=>	38700,
		30870	=>	38697,
		30871	=>	38694,
		30872	=>	38691,
		30873	=>	38688,
		30874	=>	38685,
		30875	=>	38682,
		30876	=>	38679,
		30877	=>	38676,
		30878	=>	38673,
		30879	=>	38669,
		30880	=>	38666,
		30881	=>	38663,
		30882	=>	38660,
		30883	=>	38657,
		30884	=>	38654,
		30885	=>	38651,
		30886	=>	38648,
		30887	=>	38645,
		30888	=>	38642,
		30889	=>	38639,
		30890	=>	38635,
		30891	=>	38632,
		30892	=>	38629,
		30893	=>	38626,
		30894	=>	38623,
		30895	=>	38620,
		30896	=>	38617,
		30897	=>	38614,
		30898	=>	38611,
		30899	=>	38608,
		30900	=>	38605,
		30901	=>	38601,
		30902	=>	38598,
		30903	=>	38595,
		30904	=>	38592,
		30905	=>	38589,
		30906	=>	38586,
		30907	=>	38583,
		30908	=>	38580,
		30909	=>	38577,
		30910	=>	38574,
		30911	=>	38571,
		30912	=>	38567,
		30913	=>	38564,
		30914	=>	38561,
		30915	=>	38558,
		30916	=>	38555,
		30917	=>	38552,
		30918	=>	38549,
		30919	=>	38546,
		30920	=>	38543,
		30921	=>	38540,
		30922	=>	38537,
		30923	=>	38533,
		30924	=>	38530,
		30925	=>	38527,
		30926	=>	38524,
		30927	=>	38521,
		30928	=>	38518,
		30929	=>	38515,
		30930	=>	38512,
		30931	=>	38509,
		30932	=>	38506,
		30933	=>	38503,
		30934	=>	38499,
		30935	=>	38496,
		30936	=>	38493,
		30937	=>	38490,
		30938	=>	38487,
		30939	=>	38484,
		30940	=>	38481,
		30941	=>	38478,
		30942	=>	38475,
		30943	=>	38472,
		30944	=>	38469,
		30945	=>	38465,
		30946	=>	38462,
		30947	=>	38459,
		30948	=>	38456,
		30949	=>	38453,
		30950	=>	38450,
		30951	=>	38447,
		30952	=>	38444,
		30953	=>	38441,
		30954	=>	38438,
		30955	=>	38434,
		30956	=>	38431,
		30957	=>	38428,
		30958	=>	38425,
		30959	=>	38422,
		30960	=>	38419,
		30961	=>	38416,
		30962	=>	38413,
		30963	=>	38410,
		30964	=>	38407,
		30965	=>	38404,
		30966	=>	38400,
		30967	=>	38397,
		30968	=>	38394,
		30969	=>	38391,
		30970	=>	38388,
		30971	=>	38385,
		30972	=>	38382,
		30973	=>	38379,
		30974	=>	38376,
		30975	=>	38373,
		30976	=>	38369,
		30977	=>	38366,
		30978	=>	38363,
		30979	=>	38360,
		30980	=>	38357,
		30981	=>	38354,
		30982	=>	38351,
		30983	=>	38348,
		30984	=>	38345,
		30985	=>	38342,
		30986	=>	38339,
		30987	=>	38335,
		30988	=>	38332,
		30989	=>	38329,
		30990	=>	38326,
		30991	=>	38323,
		30992	=>	38320,
		30993	=>	38317,
		30994	=>	38314,
		30995	=>	38311,
		30996	=>	38308,
		30997	=>	38304,
		30998	=>	38301,
		30999	=>	38298,
		31000	=>	38295,
		31001	=>	38292,
		31002	=>	38289,
		31003	=>	38286,
		31004	=>	38283,
		31005	=>	38280,
		31006	=>	38277,
		31007	=>	38274,
		31008	=>	38270,
		31009	=>	38267,
		31010	=>	38264,
		31011	=>	38261,
		31012	=>	38258,
		31013	=>	38255,
		31014	=>	38252,
		31015	=>	38249,
		31016	=>	38246,
		31017	=>	38243,
		31018	=>	38239,
		31019	=>	38236,
		31020	=>	38233,
		31021	=>	38230,
		31022	=>	38227,
		31023	=>	38224,
		31024	=>	38221,
		31025	=>	38218,
		31026	=>	38215,
		31027	=>	38212,
		31028	=>	38208,
		31029	=>	38205,
		31030	=>	38202,
		31031	=>	38199,
		31032	=>	38196,
		31033	=>	38193,
		31034	=>	38190,
		31035	=>	38187,
		31036	=>	38184,
		31037	=>	38181,
		31038	=>	38177,
		31039	=>	38174,
		31040	=>	38171,
		31041	=>	38168,
		31042	=>	38165,
		31043	=>	38162,
		31044	=>	38159,
		31045	=>	38156,
		31046	=>	38153,
		31047	=>	38150,
		31048	=>	38147,
		31049	=>	38143,
		31050	=>	38140,
		31051	=>	38137,
		31052	=>	38134,
		31053	=>	38131,
		31054	=>	38128,
		31055	=>	38125,
		31056	=>	38122,
		31057	=>	38119,
		31058	=>	38116,
		31059	=>	38112,
		31060	=>	38109,
		31061	=>	38106,
		31062	=>	38103,
		31063	=>	38100,
		31064	=>	38097,
		31065	=>	38094,
		31066	=>	38091,
		31067	=>	38088,
		31068	=>	38085,
		31069	=>	38081,
		31070	=>	38078,
		31071	=>	38075,
		31072	=>	38072,
		31073	=>	38069,
		31074	=>	38066,
		31075	=>	38063,
		31076	=>	38060,
		31077	=>	38057,
		31078	=>	38054,
		31079	=>	38050,
		31080	=>	38047,
		31081	=>	38044,
		31082	=>	38041,
		31083	=>	38038,
		31084	=>	38035,
		31085	=>	38032,
		31086	=>	38029,
		31087	=>	38026,
		31088	=>	38023,
		31089	=>	38019,
		31090	=>	38016,
		31091	=>	38013,
		31092	=>	38010,
		31093	=>	38007,
		31094	=>	38004,
		31095	=>	38001,
		31096	=>	37998,
		31097	=>	37995,
		31098	=>	37991,
		31099	=>	37988,
		31100	=>	37985,
		31101	=>	37982,
		31102	=>	37979,
		31103	=>	37976,
		31104	=>	37973,
		31105	=>	37970,
		31106	=>	37967,
		31107	=>	37964,
		31108	=>	37960,
		31109	=>	37957,
		31110	=>	37954,
		31111	=>	37951,
		31112	=>	37948,
		31113	=>	37945,
		31114	=>	37942,
		31115	=>	37939,
		31116	=>	37936,
		31117	=>	37933,
		31118	=>	37929,
		31119	=>	37926,
		31120	=>	37923,
		31121	=>	37920,
		31122	=>	37917,
		31123	=>	37914,
		31124	=>	37911,
		31125	=>	37908,
		31126	=>	37905,
		31127	=>	37902,
		31128	=>	37898,
		31129	=>	37895,
		31130	=>	37892,
		31131	=>	37889,
		31132	=>	37886,
		31133	=>	37883,
		31134	=>	37880,
		31135	=>	37877,
		31136	=>	37874,
		31137	=>	37871,
		31138	=>	37867,
		31139	=>	37864,
		31140	=>	37861,
		31141	=>	37858,
		31142	=>	37855,
		31143	=>	37852,
		31144	=>	37849,
		31145	=>	37846,
		31146	=>	37843,
		31147	=>	37839,
		31148	=>	37836,
		31149	=>	37833,
		31150	=>	37830,
		31151	=>	37827,
		31152	=>	37824,
		31153	=>	37821,
		31154	=>	37818,
		31155	=>	37815,
		31156	=>	37812,
		31157	=>	37808,
		31158	=>	37805,
		31159	=>	37802,
		31160	=>	37799,
		31161	=>	37796,
		31162	=>	37793,
		31163	=>	37790,
		31164	=>	37787,
		31165	=>	37784,
		31166	=>	37780,
		31167	=>	37777,
		31168	=>	37774,
		31169	=>	37771,
		31170	=>	37768,
		31171	=>	37765,
		31172	=>	37762,
		31173	=>	37759,
		31174	=>	37756,
		31175	=>	37753,
		31176	=>	37749,
		31177	=>	37746,
		31178	=>	37743,
		31179	=>	37740,
		31180	=>	37737,
		31181	=>	37734,
		31182	=>	37731,
		31183	=>	37728,
		31184	=>	37725,
		31185	=>	37721,
		31186	=>	37718,
		31187	=>	37715,
		31188	=>	37712,
		31189	=>	37709,
		31190	=>	37706,
		31191	=>	37703,
		31192	=>	37700,
		31193	=>	37697,
		31194	=>	37694,
		31195	=>	37690,
		31196	=>	37687,
		31197	=>	37684,
		31198	=>	37681,
		31199	=>	37678,
		31200	=>	37675,
		31201	=>	37672,
		31202	=>	37669,
		31203	=>	37666,
		31204	=>	37662,
		31205	=>	37659,
		31206	=>	37656,
		31207	=>	37653,
		31208	=>	37650,
		31209	=>	37647,
		31210	=>	37644,
		31211	=>	37641,
		31212	=>	37638,
		31213	=>	37635,
		31214	=>	37631,
		31215	=>	37628,
		31216	=>	37625,
		31217	=>	37622,
		31218	=>	37619,
		31219	=>	37616,
		31220	=>	37613,
		31221	=>	37610,
		31222	=>	37607,
		31223	=>	37603,
		31224	=>	37600,
		31225	=>	37597,
		31226	=>	37594,
		31227	=>	37591,
		31228	=>	37588,
		31229	=>	37585,
		31230	=>	37582,
		31231	=>	37579,
		31232	=>	37575,
		31233	=>	37572,
		31234	=>	37569,
		31235	=>	37566,
		31236	=>	37563,
		31237	=>	37560,
		31238	=>	37557,
		31239	=>	37554,
		31240	=>	37551,
		31241	=>	37548,
		31242	=>	37544,
		31243	=>	37541,
		31244	=>	37538,
		31245	=>	37535,
		31246	=>	37532,
		31247	=>	37529,
		31248	=>	37526,
		31249	=>	37523,
		31250	=>	37520,
		31251	=>	37516,
		31252	=>	37513,
		31253	=>	37510,
		31254	=>	37507,
		31255	=>	37504,
		31256	=>	37501,
		31257	=>	37498,
		31258	=>	37495,
		31259	=>	37492,
		31260	=>	37488,
		31261	=>	37485,
		31262	=>	37482,
		31263	=>	37479,
		31264	=>	37476,
		31265	=>	37473,
		31266	=>	37470,
		31267	=>	37467,
		31268	=>	37464,
		31269	=>	37460,
		31270	=>	37457,
		31271	=>	37454,
		31272	=>	37451,
		31273	=>	37448,
		31274	=>	37445,
		31275	=>	37442,
		31276	=>	37439,
		31277	=>	37436,
		31278	=>	37432,
		31279	=>	37429,
		31280	=>	37426,
		31281	=>	37423,
		31282	=>	37420,
		31283	=>	37417,
		31284	=>	37414,
		31285	=>	37411,
		31286	=>	37408,
		31287	=>	37405,
		31288	=>	37401,
		31289	=>	37398,
		31290	=>	37395,
		31291	=>	37392,
		31292	=>	37389,
		31293	=>	37386,
		31294	=>	37383,
		31295	=>	37380,
		31296	=>	37377,
		31297	=>	37373,
		31298	=>	37370,
		31299	=>	37367,
		31300	=>	37364,
		31301	=>	37361,
		31302	=>	37358,
		31303	=>	37355,
		31304	=>	37352,
		31305	=>	37349,
		31306	=>	37345,
		31307	=>	37342,
		31308	=>	37339,
		31309	=>	37336,
		31310	=>	37333,
		31311	=>	37330,
		31312	=>	37327,
		31313	=>	37324,
		31314	=>	37321,
		31315	=>	37317,
		31316	=>	37314,
		31317	=>	37311,
		31318	=>	37308,
		31319	=>	37305,
		31320	=>	37302,
		31321	=>	37299,
		31322	=>	37296,
		31323	=>	37293,
		31324	=>	37289,
		31325	=>	37286,
		31326	=>	37283,
		31327	=>	37280,
		31328	=>	37277,
		31329	=>	37274,
		31330	=>	37271,
		31331	=>	37268,
		31332	=>	37265,
		31333	=>	37261,
		31334	=>	37258,
		31335	=>	37255,
		31336	=>	37252,
		31337	=>	37249,
		31338	=>	37246,
		31339	=>	37243,
		31340	=>	37240,
		31341	=>	37237,
		31342	=>	37233,
		31343	=>	37230,
		31344	=>	37227,
		31345	=>	37224,
		31346	=>	37221,
		31347	=>	37218,
		31348	=>	37215,
		31349	=>	37212,
		31350	=>	37209,
		31351	=>	37205,
		31352	=>	37202,
		31353	=>	37199,
		31354	=>	37196,
		31355	=>	37193,
		31356	=>	37190,
		31357	=>	37187,
		31358	=>	37184,
		31359	=>	37180,
		31360	=>	37177,
		31361	=>	37174,
		31362	=>	37171,
		31363	=>	37168,
		31364	=>	37165,
		31365	=>	37162,
		31366	=>	37159,
		31367	=>	37156,
		31368	=>	37152,
		31369	=>	37149,
		31370	=>	37146,
		31371	=>	37143,
		31372	=>	37140,
		31373	=>	37137,
		31374	=>	37134,
		31375	=>	37131,
		31376	=>	37128,
		31377	=>	37124,
		31378	=>	37121,
		31379	=>	37118,
		31380	=>	37115,
		31381	=>	37112,
		31382	=>	37109,
		31383	=>	37106,
		31384	=>	37103,
		31385	=>	37100,
		31386	=>	37096,
		31387	=>	37093,
		31388	=>	37090,
		31389	=>	37087,
		31390	=>	37084,
		31391	=>	37081,
		31392	=>	37078,
		31393	=>	37075,
		31394	=>	37072,
		31395	=>	37068,
		31396	=>	37065,
		31397	=>	37062,
		31398	=>	37059,
		31399	=>	37056,
		31400	=>	37053,
		31401	=>	37050,
		31402	=>	37047,
		31403	=>	37043,
		31404	=>	37040,
		31405	=>	37037,
		31406	=>	37034,
		31407	=>	37031,
		31408	=>	37028,
		31409	=>	37025,
		31410	=>	37022,
		31411	=>	37019,
		31412	=>	37015,
		31413	=>	37012,
		31414	=>	37009,
		31415	=>	37006,
		31416	=>	37003,
		31417	=>	37000,
		31418	=>	36997,
		31419	=>	36994,
		31420	=>	36991,
		31421	=>	36987,
		31422	=>	36984,
		31423	=>	36981,
		31424	=>	36978,
		31425	=>	36975,
		31426	=>	36972,
		31427	=>	36969,
		31428	=>	36966,
		31429	=>	36962,
		31430	=>	36959,
		31431	=>	36956,
		31432	=>	36953,
		31433	=>	36950,
		31434	=>	36947,
		31435	=>	36944,
		31436	=>	36941,
		31437	=>	36938,
		31438	=>	36934,
		31439	=>	36931,
		31440	=>	36928,
		31441	=>	36925,
		31442	=>	36922,
		31443	=>	36919,
		31444	=>	36916,
		31445	=>	36913,
		31446	=>	36910,
		31447	=>	36906,
		31448	=>	36903,
		31449	=>	36900,
		31450	=>	36897,
		31451	=>	36894,
		31452	=>	36891,
		31453	=>	36888,
		31454	=>	36885,
		31455	=>	36881,
		31456	=>	36878,
		31457	=>	36875,
		31458	=>	36872,
		31459	=>	36869,
		31460	=>	36866,
		31461	=>	36863,
		31462	=>	36860,
		31463	=>	36857,
		31464	=>	36853,
		31465	=>	36850,
		31466	=>	36847,
		31467	=>	36844,
		31468	=>	36841,
		31469	=>	36838,
		31470	=>	36835,
		31471	=>	36832,
		31472	=>	36828,
		31473	=>	36825,
		31474	=>	36822,
		31475	=>	36819,
		31476	=>	36816,
		31477	=>	36813,
		31478	=>	36810,
		31479	=>	36807,
		31480	=>	36804,
		31481	=>	36800,
		31482	=>	36797,
		31483	=>	36794,
		31484	=>	36791,
		31485	=>	36788,
		31486	=>	36785,
		31487	=>	36782,
		31488	=>	36779,
		31489	=>	36775,
		31490	=>	36772,
		31491	=>	36769,
		31492	=>	36766,
		31493	=>	36763,
		31494	=>	36760,
		31495	=>	36757,
		31496	=>	36754,
		31497	=>	36751,
		31498	=>	36747,
		31499	=>	36744,
		31500	=>	36741,
		31501	=>	36738,
		31502	=>	36735,
		31503	=>	36732,
		31504	=>	36729,
		31505	=>	36726,
		31506	=>	36722,
		31507	=>	36719,
		31508	=>	36716,
		31509	=>	36713,
		31510	=>	36710,
		31511	=>	36707,
		31512	=>	36704,
		31513	=>	36701,
		31514	=>	36698,
		31515	=>	36694,
		31516	=>	36691,
		31517	=>	36688,
		31518	=>	36685,
		31519	=>	36682,
		31520	=>	36679,
		31521	=>	36676,
		31522	=>	36673,
		31523	=>	36669,
		31524	=>	36666,
		31525	=>	36663,
		31526	=>	36660,
		31527	=>	36657,
		31528	=>	36654,
		31529	=>	36651,
		31530	=>	36648,
		31531	=>	36644,
		31532	=>	36641,
		31533	=>	36638,
		31534	=>	36635,
		31535	=>	36632,
		31536	=>	36629,
		31537	=>	36626,
		31538	=>	36623,
		31539	=>	36620,
		31540	=>	36616,
		31541	=>	36613,
		31542	=>	36610,
		31543	=>	36607,
		31544	=>	36604,
		31545	=>	36601,
		31546	=>	36598,
		31547	=>	36595,
		31548	=>	36591,
		31549	=>	36588,
		31550	=>	36585,
		31551	=>	36582,
		31552	=>	36579,
		31553	=>	36576,
		31554	=>	36573,
		31555	=>	36570,
		31556	=>	36566,
		31557	=>	36563,
		31558	=>	36560,
		31559	=>	36557,
		31560	=>	36554,
		31561	=>	36551,
		31562	=>	36548,
		31563	=>	36545,
		31564	=>	36542,
		31565	=>	36538,
		31566	=>	36535,
		31567	=>	36532,
		31568	=>	36529,
		31569	=>	36526,
		31570	=>	36523,
		31571	=>	36520,
		31572	=>	36517,
		31573	=>	36513,
		31574	=>	36510,
		31575	=>	36507,
		31576	=>	36504,
		31577	=>	36501,
		31578	=>	36498,
		31579	=>	36495,
		31580	=>	36492,
		31581	=>	36488,
		31582	=>	36485,
		31583	=>	36482,
		31584	=>	36479,
		31585	=>	36476,
		31586	=>	36473,
		31587	=>	36470,
		31588	=>	36467,
		31589	=>	36463,
		31590	=>	36460,
		31591	=>	36457,
		31592	=>	36454,
		31593	=>	36451,
		31594	=>	36448,
		31595	=>	36445,
		31596	=>	36442,
		31597	=>	36439,
		31598	=>	36435,
		31599	=>	36432,
		31600	=>	36429,
		31601	=>	36426,
		31602	=>	36423,
		31603	=>	36420,
		31604	=>	36417,
		31605	=>	36414,
		31606	=>	36410,
		31607	=>	36407,
		31608	=>	36404,
		31609	=>	36401,
		31610	=>	36398,
		31611	=>	36395,
		31612	=>	36392,
		31613	=>	36389,
		31614	=>	36385,
		31615	=>	36382,
		31616	=>	36379,
		31617	=>	36376,
		31618	=>	36373,
		31619	=>	36370,
		31620	=>	36367,
		31621	=>	36364,
		31622	=>	36360,
		31623	=>	36357,
		31624	=>	36354,
		31625	=>	36351,
		31626	=>	36348,
		31627	=>	36345,
		31628	=>	36342,
		31629	=>	36339,
		31630	=>	36335,
		31631	=>	36332,
		31632	=>	36329,
		31633	=>	36326,
		31634	=>	36323,
		31635	=>	36320,
		31636	=>	36317,
		31637	=>	36314,
		31638	=>	36311,
		31639	=>	36307,
		31640	=>	36304,
		31641	=>	36301,
		31642	=>	36298,
		31643	=>	36295,
		31644	=>	36292,
		31645	=>	36289,
		31646	=>	36286,
		31647	=>	36282,
		31648	=>	36279,
		31649	=>	36276,
		31650	=>	36273,
		31651	=>	36270,
		31652	=>	36267,
		31653	=>	36264,
		31654	=>	36261,
		31655	=>	36257,
		31656	=>	36254,
		31657	=>	36251,
		31658	=>	36248,
		31659	=>	36245,
		31660	=>	36242,
		31661	=>	36239,
		31662	=>	36236,
		31663	=>	36232,
		31664	=>	36229,
		31665	=>	36226,
		31666	=>	36223,
		31667	=>	36220,
		31668	=>	36217,
		31669	=>	36214,
		31670	=>	36211,
		31671	=>	36207,
		31672	=>	36204,
		31673	=>	36201,
		31674	=>	36198,
		31675	=>	36195,
		31676	=>	36192,
		31677	=>	36189,
		31678	=>	36186,
		31679	=>	36182,
		31680	=>	36179,
		31681	=>	36176,
		31682	=>	36173,
		31683	=>	36170,
		31684	=>	36167,
		31685	=>	36164,
		31686	=>	36161,
		31687	=>	36157,
		31688	=>	36154,
		31689	=>	36151,
		31690	=>	36148,
		31691	=>	36145,
		31692	=>	36142,
		31693	=>	36139,
		31694	=>	36136,
		31695	=>	36132,
		31696	=>	36129,
		31697	=>	36126,
		31698	=>	36123,
		31699	=>	36120,
		31700	=>	36117,
		31701	=>	36114,
		31702	=>	36111,
		31703	=>	36107,
		31704	=>	36104,
		31705	=>	36101,
		31706	=>	36098,
		31707	=>	36095,
		31708	=>	36092,
		31709	=>	36089,
		31710	=>	36086,
		31711	=>	36082,
		31712	=>	36079,
		31713	=>	36076,
		31714	=>	36073,
		31715	=>	36070,
		31716	=>	36067,
		31717	=>	36064,
		31718	=>	36061,
		31719	=>	36057,
		31720	=>	36054,
		31721	=>	36051,
		31722	=>	36048,
		31723	=>	36045,
		31724	=>	36042,
		31725	=>	36039,
		31726	=>	36036,
		31727	=>	36032,
		31728	=>	36029,
		31729	=>	36026,
		31730	=>	36023,
		31731	=>	36020,
		31732	=>	36017,
		31733	=>	36014,
		31734	=>	36011,
		31735	=>	36007,
		31736	=>	36004,
		31737	=>	36001,
		31738	=>	35998,
		31739	=>	35995,
		31740	=>	35992,
		31741	=>	35989,
		31742	=>	35986,
		31743	=>	35982,
		31744	=>	35979,
		31745	=>	35976,
		31746	=>	35973,
		31747	=>	35970,
		31748	=>	35967,
		31749	=>	35964,
		31750	=>	35961,
		31751	=>	35957,
		31752	=>	35954,
		31753	=>	35951,
		31754	=>	35948,
		31755	=>	35945,
		31756	=>	35942,
		31757	=>	35939,
		31758	=>	35936,
		31759	=>	35932,
		31760	=>	35929,
		31761	=>	35926,
		31762	=>	35923,
		31763	=>	35920,
		31764	=>	35917,
		31765	=>	35914,
		31766	=>	35910,
		31767	=>	35907,
		31768	=>	35904,
		31769	=>	35901,
		31770	=>	35898,
		31771	=>	35895,
		31772	=>	35892,
		31773	=>	35889,
		31774	=>	35885,
		31775	=>	35882,
		31776	=>	35879,
		31777	=>	35876,
		31778	=>	35873,
		31779	=>	35870,
		31780	=>	35867,
		31781	=>	35864,
		31782	=>	35860,
		31783	=>	35857,
		31784	=>	35854,
		31785	=>	35851,
		31786	=>	35848,
		31787	=>	35845,
		31788	=>	35842,
		31789	=>	35839,
		31790	=>	35835,
		31791	=>	35832,
		31792	=>	35829,
		31793	=>	35826,
		31794	=>	35823,
		31795	=>	35820,
		31796	=>	35817,
		31797	=>	35814,
		31798	=>	35810,
		31799	=>	35807,
		31800	=>	35804,
		31801	=>	35801,
		31802	=>	35798,
		31803	=>	35795,
		31804	=>	35792,
		31805	=>	35789,
		31806	=>	35785,
		31807	=>	35782,
		31808	=>	35779,
		31809	=>	35776,
		31810	=>	35773,
		31811	=>	35770,
		31812	=>	35767,
		31813	=>	35763,
		31814	=>	35760,
		31815	=>	35757,
		31816	=>	35754,
		31817	=>	35751,
		31818	=>	35748,
		31819	=>	35745,
		31820	=>	35742,
		31821	=>	35738,
		31822	=>	35735,
		31823	=>	35732,
		31824	=>	35729,
		31825	=>	35726,
		31826	=>	35723,
		31827	=>	35720,
		31828	=>	35717,
		31829	=>	35713,
		31830	=>	35710,
		31831	=>	35707,
		31832	=>	35704,
		31833	=>	35701,
		31834	=>	35698,
		31835	=>	35695,
		31836	=>	35692,
		31837	=>	35688,
		31838	=>	35685,
		31839	=>	35682,
		31840	=>	35679,
		31841	=>	35676,
		31842	=>	35673,
		31843	=>	35670,
		31844	=>	35666,
		31845	=>	35663,
		31846	=>	35660,
		31847	=>	35657,
		31848	=>	35654,
		31849	=>	35651,
		31850	=>	35648,
		31851	=>	35645,
		31852	=>	35641,
		31853	=>	35638,
		31854	=>	35635,
		31855	=>	35632,
		31856	=>	35629,
		31857	=>	35626,
		31858	=>	35623,
		31859	=>	35620,
		31860	=>	35616,
		31861	=>	35613,
		31862	=>	35610,
		31863	=>	35607,
		31864	=>	35604,
		31865	=>	35601,
		31866	=>	35598,
		31867	=>	35595,
		31868	=>	35591,
		31869	=>	35588,
		31870	=>	35585,
		31871	=>	35582,
		31872	=>	35579,
		31873	=>	35576,
		31874	=>	35573,
		31875	=>	35569,
		31876	=>	35566,
		31877	=>	35563,
		31878	=>	35560,
		31879	=>	35557,
		31880	=>	35554,
		31881	=>	35551,
		31882	=>	35548,
		31883	=>	35544,
		31884	=>	35541,
		31885	=>	35538,
		31886	=>	35535,
		31887	=>	35532,
		31888	=>	35529,
		31889	=>	35526,
		31890	=>	35523,
		31891	=>	35519,
		31892	=>	35516,
		31893	=>	35513,
		31894	=>	35510,
		31895	=>	35507,
		31896	=>	35504,
		31897	=>	35501,
		31898	=>	35497,
		31899	=>	35494,
		31900	=>	35491,
		31901	=>	35488,
		31902	=>	35485,
		31903	=>	35482,
		31904	=>	35479,
		31905	=>	35476,
		31906	=>	35472,
		31907	=>	35469,
		31908	=>	35466,
		31909	=>	35463,
		31910	=>	35460,
		31911	=>	35457,
		31912	=>	35454,
		31913	=>	35451,
		31914	=>	35447,
		31915	=>	35444,
		31916	=>	35441,
		31917	=>	35438,
		31918	=>	35435,
		31919	=>	35432,
		31920	=>	35429,
		31921	=>	35425,
		31922	=>	35422,
		31923	=>	35419,
		31924	=>	35416,
		31925	=>	35413,
		31926	=>	35410,
		31927	=>	35407,
		31928	=>	35404,
		31929	=>	35400,
		31930	=>	35397,
		31931	=>	35394,
		31932	=>	35391,
		31933	=>	35388,
		31934	=>	35385,
		31935	=>	35382,
		31936	=>	35378,
		31937	=>	35375,
		31938	=>	35372,
		31939	=>	35369,
		31940	=>	35366,
		31941	=>	35363,
		31942	=>	35360,
		31943	=>	35357,
		31944	=>	35353,
		31945	=>	35350,
		31946	=>	35347,
		31947	=>	35344,
		31948	=>	35341,
		31949	=>	35338,
		31950	=>	35335,
		31951	=>	35332,
		31952	=>	35328,
		31953	=>	35325,
		31954	=>	35322,
		31955	=>	35319,
		31956	=>	35316,
		31957	=>	35313,
		31958	=>	35310,
		31959	=>	35306,
		31960	=>	35303,
		31961	=>	35300,
		31962	=>	35297,
		31963	=>	35294,
		31964	=>	35291,
		31965	=>	35288,
		31966	=>	35285,
		31967	=>	35281,
		31968	=>	35278,
		31969	=>	35275,
		31970	=>	35272,
		31971	=>	35269,
		31972	=>	35266,
		31973	=>	35263,
		31974	=>	35259,
		31975	=>	35256,
		31976	=>	35253,
		31977	=>	35250,
		31978	=>	35247,
		31979	=>	35244,
		31980	=>	35241,
		31981	=>	35238,
		31982	=>	35234,
		31983	=>	35231,
		31984	=>	35228,
		31985	=>	35225,
		31986	=>	35222,
		31987	=>	35219,
		31988	=>	35216,
		31989	=>	35212,
		31990	=>	35209,
		31991	=>	35206,
		31992	=>	35203,
		31993	=>	35200,
		31994	=>	35197,
		31995	=>	35194,
		31996	=>	35191,
		31997	=>	35187,
		31998	=>	35184,
		31999	=>	35181,
		32000	=>	35178,
		32001	=>	35175,
		32002	=>	35172,
		32003	=>	35169,
		32004	=>	35165,
		32005	=>	35162,
		32006	=>	35159,
		32007	=>	35156,
		32008	=>	35153,
		32009	=>	35150,
		32010	=>	35147,
		32011	=>	35144,
		32012	=>	35140,
		32013	=>	35137,
		32014	=>	35134,
		32015	=>	35131,
		32016	=>	35128,
		32017	=>	35125,
		32018	=>	35122,
		32019	=>	35118,
		32020	=>	35115,
		32021	=>	35112,
		32022	=>	35109,
		32023	=>	35106,
		32024	=>	35103,
		32025	=>	35100,
		32026	=>	35097,
		32027	=>	35093,
		32028	=>	35090,
		32029	=>	35087,
		32030	=>	35084,
		32031	=>	35081,
		32032	=>	35078,
		32033	=>	35075,
		32034	=>	35071,
		32035	=>	35068,
		32036	=>	35065,
		32037	=>	35062,
		32038	=>	35059,
		32039	=>	35056,
		32040	=>	35053,
		32041	=>	35050,
		32042	=>	35046,
		32043	=>	35043,
		32044	=>	35040,
		32045	=>	35037,
		32046	=>	35034,
		32047	=>	35031,
		32048	=>	35028,
		32049	=>	35024,
		32050	=>	35021,
		32051	=>	35018,
		32052	=>	35015,
		32053	=>	35012,
		32054	=>	35009,
		32055	=>	35006,
		32056	=>	35003,
		32057	=>	34999,
		32058	=>	34996,
		32059	=>	34993,
		32060	=>	34990,
		32061	=>	34987,
		32062	=>	34984,
		32063	=>	34981,
		32064	=>	34977,
		32065	=>	34974,
		32066	=>	34971,
		32067	=>	34968,
		32068	=>	34965,
		32069	=>	34962,
		32070	=>	34959,
		32071	=>	34956,
		32072	=>	34952,
		32073	=>	34949,
		32074	=>	34946,
		32075	=>	34943,
		32076	=>	34940,
		32077	=>	34937,
		32078	=>	34934,
		32079	=>	34930,
		32080	=>	34927,
		32081	=>	34924,
		32082	=>	34921,
		32083	=>	34918,
		32084	=>	34915,
		32085	=>	34912,
		32086	=>	34909,
		32087	=>	34905,
		32088	=>	34902,
		32089	=>	34899,
		32090	=>	34896,
		32091	=>	34893,
		32092	=>	34890,
		32093	=>	34887,
		32094	=>	34883,
		32095	=>	34880,
		32096	=>	34877,
		32097	=>	34874,
		32098	=>	34871,
		32099	=>	34868,
		32100	=>	34865,
		32101	=>	34861,
		32102	=>	34858,
		32103	=>	34855,
		32104	=>	34852,
		32105	=>	34849,
		32106	=>	34846,
		32107	=>	34843,
		32108	=>	34840,
		32109	=>	34836,
		32110	=>	34833,
		32111	=>	34830,
		32112	=>	34827,
		32113	=>	34824,
		32114	=>	34821,
		32115	=>	34818,
		32116	=>	34814,
		32117	=>	34811,
		32118	=>	34808,
		32119	=>	34805,
		32120	=>	34802,
		32121	=>	34799,
		32122	=>	34796,
		32123	=>	34793,
		32124	=>	34789,
		32125	=>	34786,
		32126	=>	34783,
		32127	=>	34780,
		32128	=>	34777,
		32129	=>	34774,
		32130	=>	34771,
		32131	=>	34767,
		32132	=>	34764,
		32133	=>	34761,
		32134	=>	34758,
		32135	=>	34755,
		32136	=>	34752,
		32137	=>	34749,
		32138	=>	34745,
		32139	=>	34742,
		32140	=>	34739,
		32141	=>	34736,
		32142	=>	34733,
		32143	=>	34730,
		32144	=>	34727,
		32145	=>	34724,
		32146	=>	34720,
		32147	=>	34717,
		32148	=>	34714,
		32149	=>	34711,
		32150	=>	34708,
		32151	=>	34705,
		32152	=>	34702,
		32153	=>	34698,
		32154	=>	34695,
		32155	=>	34692,
		32156	=>	34689,
		32157	=>	34686,
		32158	=>	34683,
		32159	=>	34680,
		32160	=>	34676,
		32161	=>	34673,
		32162	=>	34670,
		32163	=>	34667,
		32164	=>	34664,
		32165	=>	34661,
		32166	=>	34658,
		32167	=>	34655,
		32168	=>	34651,
		32169	=>	34648,
		32170	=>	34645,
		32171	=>	34642,
		32172	=>	34639,
		32173	=>	34636,
		32174	=>	34633,
		32175	=>	34629,
		32176	=>	34626,
		32177	=>	34623,
		32178	=>	34620,
		32179	=>	34617,
		32180	=>	34614,
		32181	=>	34611,
		32182	=>	34607,
		32183	=>	34604,
		32184	=>	34601,
		32185	=>	34598,
		32186	=>	34595,
		32187	=>	34592,
		32188	=>	34589,
		32189	=>	34586,
		32190	=>	34582,
		32191	=>	34579,
		32192	=>	34576,
		32193	=>	34573,
		32194	=>	34570,
		32195	=>	34567,
		32196	=>	34564,
		32197	=>	34560,
		32198	=>	34557,
		32199	=>	34554,
		32200	=>	34551,
		32201	=>	34548,
		32202	=>	34545,
		32203	=>	34542,
		32204	=>	34538,
		32205	=>	34535,
		32206	=>	34532,
		32207	=>	34529,
		32208	=>	34526,
		32209	=>	34523,
		32210	=>	34520,
		32211	=>	34517,
		32212	=>	34513,
		32213	=>	34510,
		32214	=>	34507,
		32215	=>	34504,
		32216	=>	34501,
		32217	=>	34498,
		32218	=>	34495,
		32219	=>	34491,
		32220	=>	34488,
		32221	=>	34485,
		32222	=>	34482,
		32223	=>	34479,
		32224	=>	34476,
		32225	=>	34473,
		32226	=>	34469,
		32227	=>	34466,
		32228	=>	34463,
		32229	=>	34460,
		32230	=>	34457,
		32231	=>	34454,
		32232	=>	34451,
		32233	=>	34447,
		32234	=>	34444,
		32235	=>	34441,
		32236	=>	34438,
		32237	=>	34435,
		32238	=>	34432,
		32239	=>	34429,
		32240	=>	34426,
		32241	=>	34422,
		32242	=>	34419,
		32243	=>	34416,
		32244	=>	34413,
		32245	=>	34410,
		32246	=>	34407,
		32247	=>	34404,
		32248	=>	34400,
		32249	=>	34397,
		32250	=>	34394,
		32251	=>	34391,
		32252	=>	34388,
		32253	=>	34385,
		32254	=>	34382,
		32255	=>	34378,
		32256	=>	34375,
		32257	=>	34372,
		32258	=>	34369,
		32259	=>	34366,
		32260	=>	34363,
		32261	=>	34360,
		32262	=>	34356,
		32263	=>	34353,
		32264	=>	34350,
		32265	=>	34347,
		32266	=>	34344,
		32267	=>	34341,
		32268	=>	34338,
		32269	=>	34335,
		32270	=>	34331,
		32271	=>	34328,
		32272	=>	34325,
		32273	=>	34322,
		32274	=>	34319,
		32275	=>	34316,
		32276	=>	34313,
		32277	=>	34309,
		32278	=>	34306,
		32279	=>	34303,
		32280	=>	34300,
		32281	=>	34297,
		32282	=>	34294,
		32283	=>	34291,
		32284	=>	34287,
		32285	=>	34284,
		32286	=>	34281,
		32287	=>	34278,
		32288	=>	34275,
		32289	=>	34272,
		32290	=>	34269,
		32291	=>	34265,
		32292	=>	34262,
		32293	=>	34259,
		32294	=>	34256,
		32295	=>	34253,
		32296	=>	34250,
		32297	=>	34247,
		32298	=>	34244,
		32299	=>	34240,
		32300	=>	34237,
		32301	=>	34234,
		32302	=>	34231,
		32303	=>	34228,
		32304	=>	34225,
		32305	=>	34222,
		32306	=>	34218,
		32307	=>	34215,
		32308	=>	34212,
		32309	=>	34209,
		32310	=>	34206,
		32311	=>	34203,
		32312	=>	34200,
		32313	=>	34196,
		32314	=>	34193,
		32315	=>	34190,
		32316	=>	34187,
		32317	=>	34184,
		32318	=>	34181,
		32319	=>	34178,
		32320	=>	34174,
		32321	=>	34171,
		32322	=>	34168,
		32323	=>	34165,
		32324	=>	34162,
		32325	=>	34159,
		32326	=>	34156,
		32327	=>	34153,
		32328	=>	34149,
		32329	=>	34146,
		32330	=>	34143,
		32331	=>	34140,
		32332	=>	34137,
		32333	=>	34134,
		32334	=>	34131,
		32335	=>	34127,
		32336	=>	34124,
		32337	=>	34121,
		32338	=>	34118,
		32339	=>	34115,
		32340	=>	34112,
		32341	=>	34109,
		32342	=>	34105,
		32343	=>	34102,
		32344	=>	34099,
		32345	=>	34096,
		32346	=>	34093,
		32347	=>	34090,
		32348	=>	34087,
		32349	=>	34083,
		32350	=>	34080,
		32351	=>	34077,
		32352	=>	34074,
		32353	=>	34071,
		32354	=>	34068,
		32355	=>	34065,
		32356	=>	34061,
		32357	=>	34058,
		32358	=>	34055,
		32359	=>	34052,
		32360	=>	34049,
		32361	=>	34046,
		32362	=>	34043,
		32363	=>	34040,
		32364	=>	34036,
		32365	=>	34033,
		32366	=>	34030,
		32367	=>	34027,
		32368	=>	34024,
		32369	=>	34021,
		32370	=>	34018,
		32371	=>	34014,
		32372	=>	34011,
		32373	=>	34008,
		32374	=>	34005,
		32375	=>	34002,
		32376	=>	33999,
		32377	=>	33996,
		32378	=>	33992,
		32379	=>	33989,
		32380	=>	33986,
		32381	=>	33983,
		32382	=>	33980,
		32383	=>	33977,
		32384	=>	33974,
		32385	=>	33970,
		32386	=>	33967,
		32387	=>	33964,
		32388	=>	33961,
		32389	=>	33958,
		32390	=>	33955,
		32391	=>	33952,
		32392	=>	33948,
		32393	=>	33945,
		32394	=>	33942,
		32395	=>	33939,
		32396	=>	33936,
		32397	=>	33933,
		32398	=>	33930,
		32399	=>	33926,
		32400	=>	33923,
		32401	=>	33920,
		32402	=>	33917,
		32403	=>	33914,
		32404	=>	33911,
		32405	=>	33908,
		32406	=>	33905,
		32407	=>	33901,
		32408	=>	33898,
		32409	=>	33895,
		32410	=>	33892,
		32411	=>	33889,
		32412	=>	33886,
		32413	=>	33883,
		32414	=>	33879,
		32415	=>	33876,
		32416	=>	33873,
		32417	=>	33870,
		32418	=>	33867,
		32419	=>	33864,
		32420	=>	33861,
		32421	=>	33857,
		32422	=>	33854,
		32423	=>	33851,
		32424	=>	33848,
		32425	=>	33845,
		32426	=>	33842,
		32427	=>	33839,
		32428	=>	33835,
		32429	=>	33832,
		32430	=>	33829,
		32431	=>	33826,
		32432	=>	33823,
		32433	=>	33820,
		32434	=>	33817,
		32435	=>	33813,
		32436	=>	33810,
		32437	=>	33807,
		32438	=>	33804,
		32439	=>	33801,
		32440	=>	33798,
		32441	=>	33795,
		32442	=>	33791,
		32443	=>	33788,
		32444	=>	33785,
		32445	=>	33782,
		32446	=>	33779,
		32447	=>	33776,
		32448	=>	33773,
		32449	=>	33769,
		32450	=>	33766,
		32451	=>	33763,
		32452	=>	33760,
		32453	=>	33757,
		32454	=>	33754,
		32455	=>	33751,
		32456	=>	33748,
		32457	=>	33744,
		32458	=>	33741,
		32459	=>	33738,
		32460	=>	33735,
		32461	=>	33732,
		32462	=>	33729,
		32463	=>	33726,
		32464	=>	33722,
		32465	=>	33719,
		32466	=>	33716,
		32467	=>	33713,
		32468	=>	33710,
		32469	=>	33707,
		32470	=>	33704,
		32471	=>	33700,
		32472	=>	33697,
		32473	=>	33694,
		32474	=>	33691,
		32475	=>	33688,
		32476	=>	33685,
		32477	=>	33682,
		32478	=>	33678,
		32479	=>	33675,
		32480	=>	33672,
		32481	=>	33669,
		32482	=>	33666,
		32483	=>	33663,
		32484	=>	33660,
		32485	=>	33656,
		32486	=>	33653,
		32487	=>	33650,
		32488	=>	33647,
		32489	=>	33644,
		32490	=>	33641,
		32491	=>	33638,
		32492	=>	33634,
		32493	=>	33631,
		32494	=>	33628,
		32495	=>	33625,
		32496	=>	33622,
		32497	=>	33619,
		32498	=>	33616,
		32499	=>	33612,
		32500	=>	33609,
		32501	=>	33606,
		32502	=>	33603,
		32503	=>	33600,
		32504	=>	33597,
		32505	=>	33594,
		32506	=>	33590,
		32507	=>	33587,
		32508	=>	33584,
		32509	=>	33581,
		32510	=>	33578,
		32511	=>	33575,
		32512	=>	33572,
		32513	=>	33569,
		32514	=>	33565,
		32515	=>	33562,
		32516	=>	33559,
		32517	=>	33556,
		32518	=>	33553,
		32519	=>	33550,
		32520	=>	33547,
		32521	=>	33543,
		32522	=>	33540,
		32523	=>	33537,
		32524	=>	33534,
		32525	=>	33531,
		32526	=>	33528,
		32527	=>	33525,
		32528	=>	33521,
		32529	=>	33518,
		32530	=>	33515,
		32531	=>	33512,
		32532	=>	33509,
		32533	=>	33506,
		32534	=>	33503,
		32535	=>	33499,
		32536	=>	33496,
		32537	=>	33493,
		32538	=>	33490,
		32539	=>	33487,
		32540	=>	33484,
		32541	=>	33481,
		32542	=>	33477,
		32543	=>	33474,
		32544	=>	33471,
		32545	=>	33468,
		32546	=>	33465,
		32547	=>	33462,
		32548	=>	33459,
		32549	=>	33455,
		32550	=>	33452,
		32551	=>	33449,
		32552	=>	33446,
		32553	=>	33443,
		32554	=>	33440,
		32555	=>	33437,
		32556	=>	33433,
		32557	=>	33430,
		32558	=>	33427,
		32559	=>	33424,
		32560	=>	33421,
		32561	=>	33418,
		32562	=>	33415,
		32563	=>	33411,
		32564	=>	33408,
		32565	=>	33405,
		32566	=>	33402,
		32567	=>	33399,
		32568	=>	33396,
		32569	=>	33393,
		32570	=>	33389,
		32571	=>	33386,
		32572	=>	33383,
		32573	=>	33380,
		32574	=>	33377,
		32575	=>	33374,
		32576	=>	33371,
		32577	=>	33368,
		32578	=>	33364,
		32579	=>	33361,
		32580	=>	33358,
		32581	=>	33355,
		32582	=>	33352,
		32583	=>	33349,
		32584	=>	33346,
		32585	=>	33342,
		32586	=>	33339,
		32587	=>	33336,
		32588	=>	33333,
		32589	=>	33330,
		32590	=>	33327,
		32591	=>	33324,
		32592	=>	33320,
		32593	=>	33317,
		32594	=>	33314,
		32595	=>	33311,
		32596	=>	33308,
		32597	=>	33305,
		32598	=>	33302,
		32599	=>	33298,
		32600	=>	33295,
		32601	=>	33292,
		32602	=>	33289,
		32603	=>	33286,
		32604	=>	33283,
		32605	=>	33280,
		32606	=>	33276,
		32607	=>	33273,
		32608	=>	33270,
		32609	=>	33267,
		32610	=>	33264,
		32611	=>	33261,
		32612	=>	33258,
		32613	=>	33254,
		32614	=>	33251,
		32615	=>	33248,
		32616	=>	33245,
		32617	=>	33242,
		32618	=>	33239,
		32619	=>	33236,
		32620	=>	33232,
		32621	=>	33229,
		32622	=>	33226,
		32623	=>	33223,
		32624	=>	33220,
		32625	=>	33217,
		32626	=>	33214,
		32627	=>	33210,
		32628	=>	33207,
		32629	=>	33204,
		32630	=>	33201,
		32631	=>	33198,
		32632	=>	33195,
		32633	=>	33192,
		32634	=>	33188,
		32635	=>	33185,
		32636	=>	33182,
		32637	=>	33179,
		32638	=>	33176,
		32639	=>	33173,
		32640	=>	33170,
		32641	=>	33166,
		32642	=>	33163,
		32643	=>	33160,
		32644	=>	33157,
		32645	=>	33154,
		32646	=>	33151,
		32647	=>	33148,
		32648	=>	33144,
		32649	=>	33141,
		32650	=>	33138,
		32651	=>	33135,
		32652	=>	33132,
		32653	=>	33129,
		32654	=>	33126,
		32655	=>	33122,
		32656	=>	33119,
		32657	=>	33116,
		32658	=>	33113,
		32659	=>	33110,
		32660	=>	33107,
		32661	=>	33104,
		32662	=>	33100,
		32663	=>	33097,
		32664	=>	33094,
		32665	=>	33091,
		32666	=>	33088,
		32667	=>	33085,
		32668	=>	33082,
		32669	=>	33079,
		32670	=>	33075,
		32671	=>	33072,
		32672	=>	33069,
		32673	=>	33066,
		32674	=>	33063,
		32675	=>	33060,
		32676	=>	33057,
		32677	=>	33053,
		32678	=>	33050,
		32679	=>	33047,
		32680	=>	33044,
		32681	=>	33041,
		32682	=>	33038,
		32683	=>	33035,
		32684	=>	33031,
		32685	=>	33028,
		32686	=>	33025,
		32687	=>	33022,
		32688	=>	33019,
		32689	=>	33016,
		32690	=>	33013,
		32691	=>	33009,
		32692	=>	33006,
		32693	=>	33003,
		32694	=>	33000,
		32695	=>	32997,
		32696	=>	32994,
		32697	=>	32991,
		32698	=>	32987,
		32699	=>	32984,
		32700	=>	32981,
		32701	=>	32978,
		32702	=>	32975,
		32703	=>	32972,
		32704	=>	32969,
		32705	=>	32965,
		32706	=>	32962,
		32707	=>	32959,
		32708	=>	32956,
		32709	=>	32953,
		32710	=>	32950,
		32711	=>	32947,
		32712	=>	32943,
		32713	=>	32940,
		32714	=>	32937,
		32715	=>	32934,
		32716	=>	32931,
		32717	=>	32928,
		32718	=>	32925,
		32719	=>	32921,
		32720	=>	32918,
		32721	=>	32915,
		32722	=>	32912,
		32723	=>	32909,
		32724	=>	32906,
		32725	=>	32903,
		32726	=>	32899,
		32727	=>	32896,
		32728	=>	32893,
		32729	=>	32890,
		32730	=>	32887,
		32731	=>	32884,
		32732	=>	32881,
		32733	=>	32877,
		32734	=>	32874,
		32735	=>	32871,
		32736	=>	32868,
		32737	=>	32865,
		32738	=>	32862,
		32739	=>	32859,
		32740	=>	32855,
		32741	=>	32852,
		32742	=>	32849,
		32743	=>	32846,
		32744	=>	32843,
		32745	=>	32840,
		32746	=>	32837,
		32747	=>	32833,
		32748	=>	32830,
		32749	=>	32827,
		32750	=>	32824,
		32751	=>	32821,
		32752	=>	32818,
		32753	=>	32815,
		32754	=>	32811,
		32755	=>	32808,
		32756	=>	32805,
		32757	=>	32802,
		32758	=>	32799,
		32759	=>	32796,
		32760	=>	32793,
		32761	=>	32789,
		32762	=>	32786,
		32763	=>	32783,
		32764	=>	32780,
		32765	=>	32777,
		32766	=>	32774,
		32767	=>	32771,
		32768	=>	32768,
		32769	=>	32764,
		32770	=>	32761,
		32771	=>	32758,
		32772	=>	32755,
		32773	=>	32752,
		32774	=>	32749,
		32775	=>	32746,
		32776	=>	32742,
		32777	=>	32739,
		32778	=>	32736,
		32779	=>	32733,
		32780	=>	32730,
		32781	=>	32727,
		32782	=>	32724,
		32783	=>	32720,
		32784	=>	32717,
		32785	=>	32714,
		32786	=>	32711,
		32787	=>	32708,
		32788	=>	32705,
		32789	=>	32702,
		32790	=>	32698,
		32791	=>	32695,
		32792	=>	32692,
		32793	=>	32689,
		32794	=>	32686,
		32795	=>	32683,
		32796	=>	32680,
		32797	=>	32676,
		32798	=>	32673,
		32799	=>	32670,
		32800	=>	32667,
		32801	=>	32664,
		32802	=>	32661,
		32803	=>	32658,
		32804	=>	32654,
		32805	=>	32651,
		32806	=>	32648,
		32807	=>	32645,
		32808	=>	32642,
		32809	=>	32639,
		32810	=>	32636,
		32811	=>	32632,
		32812	=>	32629,
		32813	=>	32626,
		32814	=>	32623,
		32815	=>	32620,
		32816	=>	32617,
		32817	=>	32614,
		32818	=>	32610,
		32819	=>	32607,
		32820	=>	32604,
		32821	=>	32601,
		32822	=>	32598,
		32823	=>	32595,
		32824	=>	32592,
		32825	=>	32588,
		32826	=>	32585,
		32827	=>	32582,
		32828	=>	32579,
		32829	=>	32576,
		32830	=>	32573,
		32831	=>	32570,
		32832	=>	32566,
		32833	=>	32563,
		32834	=>	32560,
		32835	=>	32557,
		32836	=>	32554,
		32837	=>	32551,
		32838	=>	32548,
		32839	=>	32544,
		32840	=>	32541,
		32841	=>	32538,
		32842	=>	32535,
		32843	=>	32532,
		32844	=>	32529,
		32845	=>	32526,
		32846	=>	32522,
		32847	=>	32519,
		32848	=>	32516,
		32849	=>	32513,
		32850	=>	32510,
		32851	=>	32507,
		32852	=>	32504,
		32853	=>	32500,
		32854	=>	32497,
		32855	=>	32494,
		32856	=>	32491,
		32857	=>	32488,
		32858	=>	32485,
		32859	=>	32482,
		32860	=>	32478,
		32861	=>	32475,
		32862	=>	32472,
		32863	=>	32469,
		32864	=>	32466,
		32865	=>	32463,
		32866	=>	32460,
		32867	=>	32456,
		32868	=>	32453,
		32869	=>	32450,
		32870	=>	32447,
		32871	=>	32444,
		32872	=>	32441,
		32873	=>	32438,
		32874	=>	32435,
		32875	=>	32431,
		32876	=>	32428,
		32877	=>	32425,
		32878	=>	32422,
		32879	=>	32419,
		32880	=>	32416,
		32881	=>	32413,
		32882	=>	32409,
		32883	=>	32406,
		32884	=>	32403,
		32885	=>	32400,
		32886	=>	32397,
		32887	=>	32394,
		32888	=>	32391,
		32889	=>	32387,
		32890	=>	32384,
		32891	=>	32381,
		32892	=>	32378,
		32893	=>	32375,
		32894	=>	32372,
		32895	=>	32369,
		32896	=>	32365,
		32897	=>	32362,
		32898	=>	32359,
		32899	=>	32356,
		32900	=>	32353,
		32901	=>	32350,
		32902	=>	32347,
		32903	=>	32343,
		32904	=>	32340,
		32905	=>	32337,
		32906	=>	32334,
		32907	=>	32331,
		32908	=>	32328,
		32909	=>	32325,
		32910	=>	32321,
		32911	=>	32318,
		32912	=>	32315,
		32913	=>	32312,
		32914	=>	32309,
		32915	=>	32306,
		32916	=>	32303,
		32917	=>	32299,
		32918	=>	32296,
		32919	=>	32293,
		32920	=>	32290,
		32921	=>	32287,
		32922	=>	32284,
		32923	=>	32281,
		32924	=>	32277,
		32925	=>	32274,
		32926	=>	32271,
		32927	=>	32268,
		32928	=>	32265,
		32929	=>	32262,
		32930	=>	32259,
		32931	=>	32255,
		32932	=>	32252,
		32933	=>	32249,
		32934	=>	32246,
		32935	=>	32243,
		32936	=>	32240,
		32937	=>	32237,
		32938	=>	32233,
		32939	=>	32230,
		32940	=>	32227,
		32941	=>	32224,
		32942	=>	32221,
		32943	=>	32218,
		32944	=>	32215,
		32945	=>	32211,
		32946	=>	32208,
		32947	=>	32205,
		32948	=>	32202,
		32949	=>	32199,
		32950	=>	32196,
		32951	=>	32193,
		32952	=>	32189,
		32953	=>	32186,
		32954	=>	32183,
		32955	=>	32180,
		32956	=>	32177,
		32957	=>	32174,
		32958	=>	32171,
		32959	=>	32167,
		32960	=>	32164,
		32961	=>	32161,
		32962	=>	32158,
		32963	=>	32155,
		32964	=>	32152,
		32965	=>	32149,
		32966	=>	32146,
		32967	=>	32142,
		32968	=>	32139,
		32969	=>	32136,
		32970	=>	32133,
		32971	=>	32130,
		32972	=>	32127,
		32973	=>	32124,
		32974	=>	32120,
		32975	=>	32117,
		32976	=>	32114,
		32977	=>	32111,
		32978	=>	32108,
		32979	=>	32105,
		32980	=>	32102,
		32981	=>	32098,
		32982	=>	32095,
		32983	=>	32092,
		32984	=>	32089,
		32985	=>	32086,
		32986	=>	32083,
		32987	=>	32080,
		32988	=>	32076,
		32989	=>	32073,
		32990	=>	32070,
		32991	=>	32067,
		32992	=>	32064,
		32993	=>	32061,
		32994	=>	32058,
		32995	=>	32054,
		32996	=>	32051,
		32997	=>	32048,
		32998	=>	32045,
		32999	=>	32042,
		33000	=>	32039,
		33001	=>	32036,
		33002	=>	32032,
		33003	=>	32029,
		33004	=>	32026,
		33005	=>	32023,
		33006	=>	32020,
		33007	=>	32017,
		33008	=>	32014,
		33009	=>	32010,
		33010	=>	32007,
		33011	=>	32004,
		33012	=>	32001,
		33013	=>	31998,
		33014	=>	31995,
		33015	=>	31992,
		33016	=>	31988,
		33017	=>	31985,
		33018	=>	31982,
		33019	=>	31979,
		33020	=>	31976,
		33021	=>	31973,
		33022	=>	31970,
		33023	=>	31966,
		33024	=>	31963,
		33025	=>	31960,
		33026	=>	31957,
		33027	=>	31954,
		33028	=>	31951,
		33029	=>	31948,
		33030	=>	31945,
		33031	=>	31941,
		33032	=>	31938,
		33033	=>	31935,
		33034	=>	31932,
		33035	=>	31929,
		33036	=>	31926,
		33037	=>	31923,
		33038	=>	31919,
		33039	=>	31916,
		33040	=>	31913,
		33041	=>	31910,
		33042	=>	31907,
		33043	=>	31904,
		33044	=>	31901,
		33045	=>	31897,
		33046	=>	31894,
		33047	=>	31891,
		33048	=>	31888,
		33049	=>	31885,
		33050	=>	31882,
		33051	=>	31879,
		33052	=>	31875,
		33053	=>	31872,
		33054	=>	31869,
		33055	=>	31866,
		33056	=>	31863,
		33057	=>	31860,
		33058	=>	31857,
		33059	=>	31853,
		33060	=>	31850,
		33061	=>	31847,
		33062	=>	31844,
		33063	=>	31841,
		33064	=>	31838,
		33065	=>	31835,
		33066	=>	31831,
		33067	=>	31828,
		33068	=>	31825,
		33069	=>	31822,
		33070	=>	31819,
		33071	=>	31816,
		33072	=>	31813,
		33073	=>	31809,
		33074	=>	31806,
		33075	=>	31803,
		33076	=>	31800,
		33077	=>	31797,
		33078	=>	31794,
		33079	=>	31791,
		33080	=>	31787,
		33081	=>	31784,
		33082	=>	31781,
		33083	=>	31778,
		33084	=>	31775,
		33085	=>	31772,
		33086	=>	31769,
		33087	=>	31766,
		33088	=>	31762,
		33089	=>	31759,
		33090	=>	31756,
		33091	=>	31753,
		33092	=>	31750,
		33093	=>	31747,
		33094	=>	31744,
		33095	=>	31740,
		33096	=>	31737,
		33097	=>	31734,
		33098	=>	31731,
		33099	=>	31728,
		33100	=>	31725,
		33101	=>	31722,
		33102	=>	31718,
		33103	=>	31715,
		33104	=>	31712,
		33105	=>	31709,
		33106	=>	31706,
		33107	=>	31703,
		33108	=>	31700,
		33109	=>	31696,
		33110	=>	31693,
		33111	=>	31690,
		33112	=>	31687,
		33113	=>	31684,
		33114	=>	31681,
		33115	=>	31678,
		33116	=>	31674,
		33117	=>	31671,
		33118	=>	31668,
		33119	=>	31665,
		33120	=>	31662,
		33121	=>	31659,
		33122	=>	31656,
		33123	=>	31652,
		33124	=>	31649,
		33125	=>	31646,
		33126	=>	31643,
		33127	=>	31640,
		33128	=>	31637,
		33129	=>	31634,
		33130	=>	31630,
		33131	=>	31627,
		33132	=>	31624,
		33133	=>	31621,
		33134	=>	31618,
		33135	=>	31615,
		33136	=>	31612,
		33137	=>	31609,
		33138	=>	31605,
		33139	=>	31602,
		33140	=>	31599,
		33141	=>	31596,
		33142	=>	31593,
		33143	=>	31590,
		33144	=>	31587,
		33145	=>	31583,
		33146	=>	31580,
		33147	=>	31577,
		33148	=>	31574,
		33149	=>	31571,
		33150	=>	31568,
		33151	=>	31565,
		33152	=>	31561,
		33153	=>	31558,
		33154	=>	31555,
		33155	=>	31552,
		33156	=>	31549,
		33157	=>	31546,
		33158	=>	31543,
		33159	=>	31539,
		33160	=>	31536,
		33161	=>	31533,
		33162	=>	31530,
		33163	=>	31527,
		33164	=>	31524,
		33165	=>	31521,
		33166	=>	31517,
		33167	=>	31514,
		33168	=>	31511,
		33169	=>	31508,
		33170	=>	31505,
		33171	=>	31502,
		33172	=>	31499,
		33173	=>	31495,
		33174	=>	31492,
		33175	=>	31489,
		33176	=>	31486,
		33177	=>	31483,
		33178	=>	31480,
		33179	=>	31477,
		33180	=>	31474,
		33181	=>	31470,
		33182	=>	31467,
		33183	=>	31464,
		33184	=>	31461,
		33185	=>	31458,
		33186	=>	31455,
		33187	=>	31452,
		33188	=>	31448,
		33189	=>	31445,
		33190	=>	31442,
		33191	=>	31439,
		33192	=>	31436,
		33193	=>	31433,
		33194	=>	31430,
		33195	=>	31426,
		33196	=>	31423,
		33197	=>	31420,
		33198	=>	31417,
		33199	=>	31414,
		33200	=>	31411,
		33201	=>	31408,
		33202	=>	31404,
		33203	=>	31401,
		33204	=>	31398,
		33205	=>	31395,
		33206	=>	31392,
		33207	=>	31389,
		33208	=>	31386,
		33209	=>	31382,
		33210	=>	31379,
		33211	=>	31376,
		33212	=>	31373,
		33213	=>	31370,
		33214	=>	31367,
		33215	=>	31364,
		33216	=>	31361,
		33217	=>	31357,
		33218	=>	31354,
		33219	=>	31351,
		33220	=>	31348,
		33221	=>	31345,
		33222	=>	31342,
		33223	=>	31339,
		33224	=>	31335,
		33225	=>	31332,
		33226	=>	31329,
		33227	=>	31326,
		33228	=>	31323,
		33229	=>	31320,
		33230	=>	31317,
		33231	=>	31313,
		33232	=>	31310,
		33233	=>	31307,
		33234	=>	31304,
		33235	=>	31301,
		33236	=>	31298,
		33237	=>	31295,
		33238	=>	31291,
		33239	=>	31288,
		33240	=>	31285,
		33241	=>	31282,
		33242	=>	31279,
		33243	=>	31276,
		33244	=>	31273,
		33245	=>	31270,
		33246	=>	31266,
		33247	=>	31263,
		33248	=>	31260,
		33249	=>	31257,
		33250	=>	31254,
		33251	=>	31251,
		33252	=>	31248,
		33253	=>	31244,
		33254	=>	31241,
		33255	=>	31238,
		33256	=>	31235,
		33257	=>	31232,
		33258	=>	31229,
		33259	=>	31226,
		33260	=>	31222,
		33261	=>	31219,
		33262	=>	31216,
		33263	=>	31213,
		33264	=>	31210,
		33265	=>	31207,
		33266	=>	31204,
		33267	=>	31200,
		33268	=>	31197,
		33269	=>	31194,
		33270	=>	31191,
		33271	=>	31188,
		33272	=>	31185,
		33273	=>	31182,
		33274	=>	31179,
		33275	=>	31175,
		33276	=>	31172,
		33277	=>	31169,
		33278	=>	31166,
		33279	=>	31163,
		33280	=>	31160,
		33281	=>	31157,
		33282	=>	31153,
		33283	=>	31150,
		33284	=>	31147,
		33285	=>	31144,
		33286	=>	31141,
		33287	=>	31138,
		33288	=>	31135,
		33289	=>	31131,
		33290	=>	31128,
		33291	=>	31125,
		33292	=>	31122,
		33293	=>	31119,
		33294	=>	31116,
		33295	=>	31113,
		33296	=>	31109,
		33297	=>	31106,
		33298	=>	31103,
		33299	=>	31100,
		33300	=>	31097,
		33301	=>	31094,
		33302	=>	31091,
		33303	=>	31088,
		33304	=>	31084,
		33305	=>	31081,
		33306	=>	31078,
		33307	=>	31075,
		33308	=>	31072,
		33309	=>	31069,
		33310	=>	31066,
		33311	=>	31062,
		33312	=>	31059,
		33313	=>	31056,
		33314	=>	31053,
		33315	=>	31050,
		33316	=>	31047,
		33317	=>	31044,
		33318	=>	31040,
		33319	=>	31037,
		33320	=>	31034,
		33321	=>	31031,
		33322	=>	31028,
		33323	=>	31025,
		33324	=>	31022,
		33325	=>	31018,
		33326	=>	31015,
		33327	=>	31012,
		33328	=>	31009,
		33329	=>	31006,
		33330	=>	31003,
		33331	=>	31000,
		33332	=>	30997,
		33333	=>	30993,
		33334	=>	30990,
		33335	=>	30987,
		33336	=>	30984,
		33337	=>	30981,
		33338	=>	30978,
		33339	=>	30975,
		33340	=>	30971,
		33341	=>	30968,
		33342	=>	30965,
		33343	=>	30962,
		33344	=>	30959,
		33345	=>	30956,
		33346	=>	30953,
		33347	=>	30949,
		33348	=>	30946,
		33349	=>	30943,
		33350	=>	30940,
		33351	=>	30937,
		33352	=>	30934,
		33353	=>	30931,
		33354	=>	30928,
		33355	=>	30924,
		33356	=>	30921,
		33357	=>	30918,
		33358	=>	30915,
		33359	=>	30912,
		33360	=>	30909,
		33361	=>	30906,
		33362	=>	30902,
		33363	=>	30899,
		33364	=>	30896,
		33365	=>	30893,
		33366	=>	30890,
		33367	=>	30887,
		33368	=>	30884,
		33369	=>	30880,
		33370	=>	30877,
		33371	=>	30874,
		33372	=>	30871,
		33373	=>	30868,
		33374	=>	30865,
		33375	=>	30862,
		33376	=>	30859,
		33377	=>	30855,
		33378	=>	30852,
		33379	=>	30849,
		33380	=>	30846,
		33381	=>	30843,
		33382	=>	30840,
		33383	=>	30837,
		33384	=>	30833,
		33385	=>	30830,
		33386	=>	30827,
		33387	=>	30824,
		33388	=>	30821,
		33389	=>	30818,
		33390	=>	30815,
		33391	=>	30811,
		33392	=>	30808,
		33393	=>	30805,
		33394	=>	30802,
		33395	=>	30799,
		33396	=>	30796,
		33397	=>	30793,
		33398	=>	30790,
		33399	=>	30786,
		33400	=>	30783,
		33401	=>	30780,
		33402	=>	30777,
		33403	=>	30774,
		33404	=>	30771,
		33405	=>	30768,
		33406	=>	30764,
		33407	=>	30761,
		33408	=>	30758,
		33409	=>	30755,
		33410	=>	30752,
		33411	=>	30749,
		33412	=>	30746,
		33413	=>	30742,
		33414	=>	30739,
		33415	=>	30736,
		33416	=>	30733,
		33417	=>	30730,
		33418	=>	30727,
		33419	=>	30724,
		33420	=>	30721,
		33421	=>	30717,
		33422	=>	30714,
		33423	=>	30711,
		33424	=>	30708,
		33425	=>	30705,
		33426	=>	30702,
		33427	=>	30699,
		33428	=>	30695,
		33429	=>	30692,
		33430	=>	30689,
		33431	=>	30686,
		33432	=>	30683,
		33433	=>	30680,
		33434	=>	30677,
		33435	=>	30674,
		33436	=>	30670,
		33437	=>	30667,
		33438	=>	30664,
		33439	=>	30661,
		33440	=>	30658,
		33441	=>	30655,
		33442	=>	30652,
		33443	=>	30648,
		33444	=>	30645,
		33445	=>	30642,
		33446	=>	30639,
		33447	=>	30636,
		33448	=>	30633,
		33449	=>	30630,
		33450	=>	30626,
		33451	=>	30623,
		33452	=>	30620,
		33453	=>	30617,
		33454	=>	30614,
		33455	=>	30611,
		33456	=>	30608,
		33457	=>	30605,
		33458	=>	30601,
		33459	=>	30598,
		33460	=>	30595,
		33461	=>	30592,
		33462	=>	30589,
		33463	=>	30586,
		33464	=>	30583,
		33465	=>	30579,
		33466	=>	30576,
		33467	=>	30573,
		33468	=>	30570,
		33469	=>	30567,
		33470	=>	30564,
		33471	=>	30561,
		33472	=>	30558,
		33473	=>	30554,
		33474	=>	30551,
		33475	=>	30548,
		33476	=>	30545,
		33477	=>	30542,
		33478	=>	30539,
		33479	=>	30536,
		33480	=>	30532,
		33481	=>	30529,
		33482	=>	30526,
		33483	=>	30523,
		33484	=>	30520,
		33485	=>	30517,
		33486	=>	30514,
		33487	=>	30511,
		33488	=>	30507,
		33489	=>	30504,
		33490	=>	30501,
		33491	=>	30498,
		33492	=>	30495,
		33493	=>	30492,
		33494	=>	30489,
		33495	=>	30485,
		33496	=>	30482,
		33497	=>	30479,
		33498	=>	30476,
		33499	=>	30473,
		33500	=>	30470,
		33501	=>	30467,
		33502	=>	30464,
		33503	=>	30460,
		33504	=>	30457,
		33505	=>	30454,
		33506	=>	30451,
		33507	=>	30448,
		33508	=>	30445,
		33509	=>	30442,
		33510	=>	30438,
		33511	=>	30435,
		33512	=>	30432,
		33513	=>	30429,
		33514	=>	30426,
		33515	=>	30423,
		33516	=>	30420,
		33517	=>	30417,
		33518	=>	30413,
		33519	=>	30410,
		33520	=>	30407,
		33521	=>	30404,
		33522	=>	30401,
		33523	=>	30398,
		33524	=>	30395,
		33525	=>	30391,
		33526	=>	30388,
		33527	=>	30385,
		33528	=>	30382,
		33529	=>	30379,
		33530	=>	30376,
		33531	=>	30373,
		33532	=>	30370,
		33533	=>	30366,
		33534	=>	30363,
		33535	=>	30360,
		33536	=>	30357,
		33537	=>	30354,
		33538	=>	30351,
		33539	=>	30348,
		33540	=>	30344,
		33541	=>	30341,
		33542	=>	30338,
		33543	=>	30335,
		33544	=>	30332,
		33545	=>	30329,
		33546	=>	30326,
		33547	=>	30323,
		33548	=>	30319,
		33549	=>	30316,
		33550	=>	30313,
		33551	=>	30310,
		33552	=>	30307,
		33553	=>	30304,
		33554	=>	30301,
		33555	=>	30297,
		33556	=>	30294,
		33557	=>	30291,
		33558	=>	30288,
		33559	=>	30285,
		33560	=>	30282,
		33561	=>	30279,
		33562	=>	30276,
		33563	=>	30272,
		33564	=>	30269,
		33565	=>	30266,
		33566	=>	30263,
		33567	=>	30260,
		33568	=>	30257,
		33569	=>	30254,
		33570	=>	30250,
		33571	=>	30247,
		33572	=>	30244,
		33573	=>	30241,
		33574	=>	30238,
		33575	=>	30235,
		33576	=>	30232,
		33577	=>	30229,
		33578	=>	30225,
		33579	=>	30222,
		33580	=>	30219,
		33581	=>	30216,
		33582	=>	30213,
		33583	=>	30210,
		33584	=>	30207,
		33585	=>	30203,
		33586	=>	30200,
		33587	=>	30197,
		33588	=>	30194,
		33589	=>	30191,
		33590	=>	30188,
		33591	=>	30185,
		33592	=>	30182,
		33593	=>	30178,
		33594	=>	30175,
		33595	=>	30172,
		33596	=>	30169,
		33597	=>	30166,
		33598	=>	30163,
		33599	=>	30160,
		33600	=>	30157,
		33601	=>	30153,
		33602	=>	30150,
		33603	=>	30147,
		33604	=>	30144,
		33605	=>	30141,
		33606	=>	30138,
		33607	=>	30135,
		33608	=>	30131,
		33609	=>	30128,
		33610	=>	30125,
		33611	=>	30122,
		33612	=>	30119,
		33613	=>	30116,
		33614	=>	30113,
		33615	=>	30110,
		33616	=>	30106,
		33617	=>	30103,
		33618	=>	30100,
		33619	=>	30097,
		33620	=>	30094,
		33621	=>	30091,
		33622	=>	30088,
		33623	=>	30084,
		33624	=>	30081,
		33625	=>	30078,
		33626	=>	30075,
		33627	=>	30072,
		33628	=>	30069,
		33629	=>	30066,
		33630	=>	30063,
		33631	=>	30059,
		33632	=>	30056,
		33633	=>	30053,
		33634	=>	30050,
		33635	=>	30047,
		33636	=>	30044,
		33637	=>	30041,
		33638	=>	30038,
		33639	=>	30034,
		33640	=>	30031,
		33641	=>	30028,
		33642	=>	30025,
		33643	=>	30022,
		33644	=>	30019,
		33645	=>	30016,
		33646	=>	30012,
		33647	=>	30009,
		33648	=>	30006,
		33649	=>	30003,
		33650	=>	30000,
		33651	=>	29997,
		33652	=>	29994,
		33653	=>	29991,
		33654	=>	29987,
		33655	=>	29984,
		33656	=>	29981,
		33657	=>	29978,
		33658	=>	29975,
		33659	=>	29972,
		33660	=>	29969,
		33661	=>	29966,
		33662	=>	29962,
		33663	=>	29959,
		33664	=>	29956,
		33665	=>	29953,
		33666	=>	29950,
		33667	=>	29947,
		33668	=>	29944,
		33669	=>	29940,
		33670	=>	29937,
		33671	=>	29934,
		33672	=>	29931,
		33673	=>	29928,
		33674	=>	29925,
		33675	=>	29922,
		33676	=>	29919,
		33677	=>	29915,
		33678	=>	29912,
		33679	=>	29909,
		33680	=>	29906,
		33681	=>	29903,
		33682	=>	29900,
		33683	=>	29897,
		33684	=>	29894,
		33685	=>	29890,
		33686	=>	29887,
		33687	=>	29884,
		33688	=>	29881,
		33689	=>	29878,
		33690	=>	29875,
		33691	=>	29872,
		33692	=>	29869,
		33693	=>	29865,
		33694	=>	29862,
		33695	=>	29859,
		33696	=>	29856,
		33697	=>	29853,
		33698	=>	29850,
		33699	=>	29847,
		33700	=>	29843,
		33701	=>	29840,
		33702	=>	29837,
		33703	=>	29834,
		33704	=>	29831,
		33705	=>	29828,
		33706	=>	29825,
		33707	=>	29822,
		33708	=>	29818,
		33709	=>	29815,
		33710	=>	29812,
		33711	=>	29809,
		33712	=>	29806,
		33713	=>	29803,
		33714	=>	29800,
		33715	=>	29797,
		33716	=>	29793,
		33717	=>	29790,
		33718	=>	29787,
		33719	=>	29784,
		33720	=>	29781,
		33721	=>	29778,
		33722	=>	29775,
		33723	=>	29772,
		33724	=>	29768,
		33725	=>	29765,
		33726	=>	29762,
		33727	=>	29759,
		33728	=>	29756,
		33729	=>	29753,
		33730	=>	29750,
		33731	=>	29746,
		33732	=>	29743,
		33733	=>	29740,
		33734	=>	29737,
		33735	=>	29734,
		33736	=>	29731,
		33737	=>	29728,
		33738	=>	29725,
		33739	=>	29721,
		33740	=>	29718,
		33741	=>	29715,
		33742	=>	29712,
		33743	=>	29709,
		33744	=>	29706,
		33745	=>	29703,
		33746	=>	29700,
		33747	=>	29696,
		33748	=>	29693,
		33749	=>	29690,
		33750	=>	29687,
		33751	=>	29684,
		33752	=>	29681,
		33753	=>	29678,
		33754	=>	29675,
		33755	=>	29671,
		33756	=>	29668,
		33757	=>	29665,
		33758	=>	29662,
		33759	=>	29659,
		33760	=>	29656,
		33761	=>	29653,
		33762	=>	29650,
		33763	=>	29646,
		33764	=>	29643,
		33765	=>	29640,
		33766	=>	29637,
		33767	=>	29634,
		33768	=>	29631,
		33769	=>	29628,
		33770	=>	29625,
		33771	=>	29621,
		33772	=>	29618,
		33773	=>	29615,
		33774	=>	29612,
		33775	=>	29609,
		33776	=>	29606,
		33777	=>	29603,
		33778	=>	29599,
		33779	=>	29596,
		33780	=>	29593,
		33781	=>	29590,
		33782	=>	29587,
		33783	=>	29584,
		33784	=>	29581,
		33785	=>	29578,
		33786	=>	29574,
		33787	=>	29571,
		33788	=>	29568,
		33789	=>	29565,
		33790	=>	29562,
		33791	=>	29559,
		33792	=>	29556,
		33793	=>	29553,
		33794	=>	29549,
		33795	=>	29546,
		33796	=>	29543,
		33797	=>	29540,
		33798	=>	29537,
		33799	=>	29534,
		33800	=>	29531,
		33801	=>	29528,
		33802	=>	29524,
		33803	=>	29521,
		33804	=>	29518,
		33805	=>	29515,
		33806	=>	29512,
		33807	=>	29509,
		33808	=>	29506,
		33809	=>	29503,
		33810	=>	29499,
		33811	=>	29496,
		33812	=>	29493,
		33813	=>	29490,
		33814	=>	29487,
		33815	=>	29484,
		33816	=>	29481,
		33817	=>	29478,
		33818	=>	29474,
		33819	=>	29471,
		33820	=>	29468,
		33821	=>	29465,
		33822	=>	29462,
		33823	=>	29459,
		33824	=>	29456,
		33825	=>	29453,
		33826	=>	29449,
		33827	=>	29446,
		33828	=>	29443,
		33829	=>	29440,
		33830	=>	29437,
		33831	=>	29434,
		33832	=>	29431,
		33833	=>	29428,
		33834	=>	29424,
		33835	=>	29421,
		33836	=>	29418,
		33837	=>	29415,
		33838	=>	29412,
		33839	=>	29409,
		33840	=>	29406,
		33841	=>	29403,
		33842	=>	29399,
		33843	=>	29396,
		33844	=>	29393,
		33845	=>	29390,
		33846	=>	29387,
		33847	=>	29384,
		33848	=>	29381,
		33849	=>	29378,
		33850	=>	29374,
		33851	=>	29371,
		33852	=>	29368,
		33853	=>	29365,
		33854	=>	29362,
		33855	=>	29359,
		33856	=>	29356,
		33857	=>	29353,
		33858	=>	29349,
		33859	=>	29346,
		33860	=>	29343,
		33861	=>	29340,
		33862	=>	29337,
		33863	=>	29334,
		33864	=>	29331,
		33865	=>	29328,
		33866	=>	29324,
		33867	=>	29321,
		33868	=>	29318,
		33869	=>	29315,
		33870	=>	29312,
		33871	=>	29309,
		33872	=>	29306,
		33873	=>	29303,
		33874	=>	29299,
		33875	=>	29296,
		33876	=>	29293,
		33877	=>	29290,
		33878	=>	29287,
		33879	=>	29284,
		33880	=>	29281,
		33881	=>	29278,
		33882	=>	29274,
		33883	=>	29271,
		33884	=>	29268,
		33885	=>	29265,
		33886	=>	29262,
		33887	=>	29259,
		33888	=>	29256,
		33889	=>	29253,
		33890	=>	29249,
		33891	=>	29246,
		33892	=>	29243,
		33893	=>	29240,
		33894	=>	29237,
		33895	=>	29234,
		33896	=>	29231,
		33897	=>	29228,
		33898	=>	29224,
		33899	=>	29221,
		33900	=>	29218,
		33901	=>	29215,
		33902	=>	29212,
		33903	=>	29209,
		33904	=>	29206,
		33905	=>	29203,
		33906	=>	29200,
		33907	=>	29196,
		33908	=>	29193,
		33909	=>	29190,
		33910	=>	29187,
		33911	=>	29184,
		33912	=>	29181,
		33913	=>	29178,
		33914	=>	29175,
		33915	=>	29171,
		33916	=>	29168,
		33917	=>	29165,
		33918	=>	29162,
		33919	=>	29159,
		33920	=>	29156,
		33921	=>	29153,
		33922	=>	29150,
		33923	=>	29146,
		33924	=>	29143,
		33925	=>	29140,
		33926	=>	29137,
		33927	=>	29134,
		33928	=>	29131,
		33929	=>	29128,
		33930	=>	29125,
		33931	=>	29121,
		33932	=>	29118,
		33933	=>	29115,
		33934	=>	29112,
		33935	=>	29109,
		33936	=>	29106,
		33937	=>	29103,
		33938	=>	29100,
		33939	=>	29096,
		33940	=>	29093,
		33941	=>	29090,
		33942	=>	29087,
		33943	=>	29084,
		33944	=>	29081,
		33945	=>	29078,
		33946	=>	29075,
		33947	=>	29072,
		33948	=>	29068,
		33949	=>	29065,
		33950	=>	29062,
		33951	=>	29059,
		33952	=>	29056,
		33953	=>	29053,
		33954	=>	29050,
		33955	=>	29047,
		33956	=>	29043,
		33957	=>	29040,
		33958	=>	29037,
		33959	=>	29034,
		33960	=>	29031,
		33961	=>	29028,
		33962	=>	29025,
		33963	=>	29022,
		33964	=>	29018,
		33965	=>	29015,
		33966	=>	29012,
		33967	=>	29009,
		33968	=>	29006,
		33969	=>	29003,
		33970	=>	29000,
		33971	=>	28997,
		33972	=>	28993,
		33973	=>	28990,
		33974	=>	28987,
		33975	=>	28984,
		33976	=>	28981,
		33977	=>	28978,
		33978	=>	28975,
		33979	=>	28972,
		33980	=>	28969,
		33981	=>	28965,
		33982	=>	28962,
		33983	=>	28959,
		33984	=>	28956,
		33985	=>	28953,
		33986	=>	28950,
		33987	=>	28947,
		33988	=>	28944,
		33989	=>	28940,
		33990	=>	28937,
		33991	=>	28934,
		33992	=>	28931,
		33993	=>	28928,
		33994	=>	28925,
		33995	=>	28922,
		33996	=>	28919,
		33997	=>	28915,
		33998	=>	28912,
		33999	=>	28909,
		34000	=>	28906,
		34001	=>	28903,
		34002	=>	28900,
		34003	=>	28897,
		34004	=>	28894,
		34005	=>	28891,
		34006	=>	28887,
		34007	=>	28884,
		34008	=>	28881,
		34009	=>	28878,
		34010	=>	28875,
		34011	=>	28872,
		34012	=>	28869,
		34013	=>	28866,
		34014	=>	28862,
		34015	=>	28859,
		34016	=>	28856,
		34017	=>	28853,
		34018	=>	28850,
		34019	=>	28847,
		34020	=>	28844,
		34021	=>	28841,
		34022	=>	28837,
		34023	=>	28834,
		34024	=>	28831,
		34025	=>	28828,
		34026	=>	28825,
		34027	=>	28822,
		34028	=>	28819,
		34029	=>	28816,
		34030	=>	28813,
		34031	=>	28809,
		34032	=>	28806,
		34033	=>	28803,
		34034	=>	28800,
		34035	=>	28797,
		34036	=>	28794,
		34037	=>	28791,
		34038	=>	28788,
		34039	=>	28784,
		34040	=>	28781,
		34041	=>	28778,
		34042	=>	28775,
		34043	=>	28772,
		34044	=>	28769,
		34045	=>	28766,
		34046	=>	28763,
		34047	=>	28760,
		34048	=>	28756,
		34049	=>	28753,
		34050	=>	28750,
		34051	=>	28747,
		34052	=>	28744,
		34053	=>	28741,
		34054	=>	28738,
		34055	=>	28735,
		34056	=>	28731,
		34057	=>	28728,
		34058	=>	28725,
		34059	=>	28722,
		34060	=>	28719,
		34061	=>	28716,
		34062	=>	28713,
		34063	=>	28710,
		34064	=>	28707,
		34065	=>	28703,
		34066	=>	28700,
		34067	=>	28697,
		34068	=>	28694,
		34069	=>	28691,
		34070	=>	28688,
		34071	=>	28685,
		34072	=>	28682,
		34073	=>	28678,
		34074	=>	28675,
		34075	=>	28672,
		34076	=>	28669,
		34077	=>	28666,
		34078	=>	28663,
		34079	=>	28660,
		34080	=>	28657,
		34081	=>	28654,
		34082	=>	28650,
		34083	=>	28647,
		34084	=>	28644,
		34085	=>	28641,
		34086	=>	28638,
		34087	=>	28635,
		34088	=>	28632,
		34089	=>	28629,
		34090	=>	28625,
		34091	=>	28622,
		34092	=>	28619,
		34093	=>	28616,
		34094	=>	28613,
		34095	=>	28610,
		34096	=>	28607,
		34097	=>	28604,
		34098	=>	28601,
		34099	=>	28597,
		34100	=>	28594,
		34101	=>	28591,
		34102	=>	28588,
		34103	=>	28585,
		34104	=>	28582,
		34105	=>	28579,
		34106	=>	28576,
		34107	=>	28573,
		34108	=>	28569,
		34109	=>	28566,
		34110	=>	28563,
		34111	=>	28560,
		34112	=>	28557,
		34113	=>	28554,
		34114	=>	28551,
		34115	=>	28548,
		34116	=>	28544,
		34117	=>	28541,
		34118	=>	28538,
		34119	=>	28535,
		34120	=>	28532,
		34121	=>	28529,
		34122	=>	28526,
		34123	=>	28523,
		34124	=>	28520,
		34125	=>	28516,
		34126	=>	28513,
		34127	=>	28510,
		34128	=>	28507,
		34129	=>	28504,
		34130	=>	28501,
		34131	=>	28498,
		34132	=>	28495,
		34133	=>	28492,
		34134	=>	28488,
		34135	=>	28485,
		34136	=>	28482,
		34137	=>	28479,
		34138	=>	28476,
		34139	=>	28473,
		34140	=>	28470,
		34141	=>	28467,
		34142	=>	28463,
		34143	=>	28460,
		34144	=>	28457,
		34145	=>	28454,
		34146	=>	28451,
		34147	=>	28448,
		34148	=>	28445,
		34149	=>	28442,
		34150	=>	28439,
		34151	=>	28435,
		34152	=>	28432,
		34153	=>	28429,
		34154	=>	28426,
		34155	=>	28423,
		34156	=>	28420,
		34157	=>	28417,
		34158	=>	28414,
		34159	=>	28411,
		34160	=>	28407,
		34161	=>	28404,
		34162	=>	28401,
		34163	=>	28398,
		34164	=>	28395,
		34165	=>	28392,
		34166	=>	28389,
		34167	=>	28386,
		34168	=>	28383,
		34169	=>	28379,
		34170	=>	28376,
		34171	=>	28373,
		34172	=>	28370,
		34173	=>	28367,
		34174	=>	28364,
		34175	=>	28361,
		34176	=>	28358,
		34177	=>	28355,
		34178	=>	28351,
		34179	=>	28348,
		34180	=>	28345,
		34181	=>	28342,
		34182	=>	28339,
		34183	=>	28336,
		34184	=>	28333,
		34185	=>	28330,
		34186	=>	28326,
		34187	=>	28323,
		34188	=>	28320,
		34189	=>	28317,
		34190	=>	28314,
		34191	=>	28311,
		34192	=>	28308,
		34193	=>	28305,
		34194	=>	28302,
		34195	=>	28298,
		34196	=>	28295,
		34197	=>	28292,
		34198	=>	28289,
		34199	=>	28286,
		34200	=>	28283,
		34201	=>	28280,
		34202	=>	28277,
		34203	=>	28274,
		34204	=>	28270,
		34205	=>	28267,
		34206	=>	28264,
		34207	=>	28261,
		34208	=>	28258,
		34209	=>	28255,
		34210	=>	28252,
		34211	=>	28249,
		34212	=>	28246,
		34213	=>	28242,
		34214	=>	28239,
		34215	=>	28236,
		34216	=>	28233,
		34217	=>	28230,
		34218	=>	28227,
		34219	=>	28224,
		34220	=>	28221,
		34221	=>	28218,
		34222	=>	28214,
		34223	=>	28211,
		34224	=>	28208,
		34225	=>	28205,
		34226	=>	28202,
		34227	=>	28199,
		34228	=>	28196,
		34229	=>	28193,
		34230	=>	28190,
		34231	=>	28186,
		34232	=>	28183,
		34233	=>	28180,
		34234	=>	28177,
		34235	=>	28174,
		34236	=>	28171,
		34237	=>	28168,
		34238	=>	28165,
		34239	=>	28162,
		34240	=>	28158,
		34241	=>	28155,
		34242	=>	28152,
		34243	=>	28149,
		34244	=>	28146,
		34245	=>	28143,
		34246	=>	28140,
		34247	=>	28137,
		34248	=>	28134,
		34249	=>	28130,
		34250	=>	28127,
		34251	=>	28124,
		34252	=>	28121,
		34253	=>	28118,
		34254	=>	28115,
		34255	=>	28112,
		34256	=>	28109,
		34257	=>	28106,
		34258	=>	28103,
		34259	=>	28099,
		34260	=>	28096,
		34261	=>	28093,
		34262	=>	28090,
		34263	=>	28087,
		34264	=>	28084,
		34265	=>	28081,
		34266	=>	28078,
		34267	=>	28075,
		34268	=>	28071,
		34269	=>	28068,
		34270	=>	28065,
		34271	=>	28062,
		34272	=>	28059,
		34273	=>	28056,
		34274	=>	28053,
		34275	=>	28050,
		34276	=>	28047,
		34277	=>	28043,
		34278	=>	28040,
		34279	=>	28037,
		34280	=>	28034,
		34281	=>	28031,
		34282	=>	28028,
		34283	=>	28025,
		34284	=>	28022,
		34285	=>	28019,
		34286	=>	28015,
		34287	=>	28012,
		34288	=>	28009,
		34289	=>	28006,
		34290	=>	28003,
		34291	=>	28000,
		34292	=>	27997,
		34293	=>	27994,
		34294	=>	27991,
		34295	=>	27987,
		34296	=>	27984,
		34297	=>	27981,
		34298	=>	27978,
		34299	=>	27975,
		34300	=>	27972,
		34301	=>	27969,
		34302	=>	27966,
		34303	=>	27963,
		34304	=>	27960,
		34305	=>	27956,
		34306	=>	27953,
		34307	=>	27950,
		34308	=>	27947,
		34309	=>	27944,
		34310	=>	27941,
		34311	=>	27938,
		34312	=>	27935,
		34313	=>	27932,
		34314	=>	27928,
		34315	=>	27925,
		34316	=>	27922,
		34317	=>	27919,
		34318	=>	27916,
		34319	=>	27913,
		34320	=>	27910,
		34321	=>	27907,
		34322	=>	27904,
		34323	=>	27900,
		34324	=>	27897,
		34325	=>	27894,
		34326	=>	27891,
		34327	=>	27888,
		34328	=>	27885,
		34329	=>	27882,
		34330	=>	27879,
		34331	=>	27876,
		34332	=>	27873,
		34333	=>	27869,
		34334	=>	27866,
		34335	=>	27863,
		34336	=>	27860,
		34337	=>	27857,
		34338	=>	27854,
		34339	=>	27851,
		34340	=>	27848,
		34341	=>	27845,
		34342	=>	27841,
		34343	=>	27838,
		34344	=>	27835,
		34345	=>	27832,
		34346	=>	27829,
		34347	=>	27826,
		34348	=>	27823,
		34349	=>	27820,
		34350	=>	27817,
		34351	=>	27814,
		34352	=>	27810,
		34353	=>	27807,
		34354	=>	27804,
		34355	=>	27801,
		34356	=>	27798,
		34357	=>	27795,
		34358	=>	27792,
		34359	=>	27789,
		34360	=>	27786,
		34361	=>	27782,
		34362	=>	27779,
		34363	=>	27776,
		34364	=>	27773,
		34365	=>	27770,
		34366	=>	27767,
		34367	=>	27764,
		34368	=>	27761,
		34369	=>	27758,
		34370	=>	27755,
		34371	=>	27751,
		34372	=>	27748,
		34373	=>	27745,
		34374	=>	27742,
		34375	=>	27739,
		34376	=>	27736,
		34377	=>	27733,
		34378	=>	27730,
		34379	=>	27727,
		34380	=>	27723,
		34381	=>	27720,
		34382	=>	27717,
		34383	=>	27714,
		34384	=>	27711,
		34385	=>	27708,
		34386	=>	27705,
		34387	=>	27702,
		34388	=>	27699,
		34389	=>	27696,
		34390	=>	27692,
		34391	=>	27689,
		34392	=>	27686,
		34393	=>	27683,
		34394	=>	27680,
		34395	=>	27677,
		34396	=>	27674,
		34397	=>	27671,
		34398	=>	27668,
		34399	=>	27664,
		34400	=>	27661,
		34401	=>	27658,
		34402	=>	27655,
		34403	=>	27652,
		34404	=>	27649,
		34405	=>	27646,
		34406	=>	27643,
		34407	=>	27640,
		34408	=>	27637,
		34409	=>	27633,
		34410	=>	27630,
		34411	=>	27627,
		34412	=>	27624,
		34413	=>	27621,
		34414	=>	27618,
		34415	=>	27615,
		34416	=>	27612,
		34417	=>	27609,
		34418	=>	27606,
		34419	=>	27602,
		34420	=>	27599,
		34421	=>	27596,
		34422	=>	27593,
		34423	=>	27590,
		34424	=>	27587,
		34425	=>	27584,
		34426	=>	27581,
		34427	=>	27578,
		34428	=>	27575,
		34429	=>	27571,
		34430	=>	27568,
		34431	=>	27565,
		34432	=>	27562,
		34433	=>	27559,
		34434	=>	27556,
		34435	=>	27553,
		34436	=>	27550,
		34437	=>	27547,
		34438	=>	27544,
		34439	=>	27540,
		34440	=>	27537,
		34441	=>	27534,
		34442	=>	27531,
		34443	=>	27528,
		34444	=>	27525,
		34445	=>	27522,
		34446	=>	27519,
		34447	=>	27516,
		34448	=>	27512,
		34449	=>	27509,
		34450	=>	27506,
		34451	=>	27503,
		34452	=>	27500,
		34453	=>	27497,
		34454	=>	27494,
		34455	=>	27491,
		34456	=>	27488,
		34457	=>	27485,
		34458	=>	27481,
		34459	=>	27478,
		34460	=>	27475,
		34461	=>	27472,
		34462	=>	27469,
		34463	=>	27466,
		34464	=>	27463,
		34465	=>	27460,
		34466	=>	27457,
		34467	=>	27454,
		34468	=>	27450,
		34469	=>	27447,
		34470	=>	27444,
		34471	=>	27441,
		34472	=>	27438,
		34473	=>	27435,
		34474	=>	27432,
		34475	=>	27429,
		34476	=>	27426,
		34477	=>	27423,
		34478	=>	27419,
		34479	=>	27416,
		34480	=>	27413,
		34481	=>	27410,
		34482	=>	27407,
		34483	=>	27404,
		34484	=>	27401,
		34485	=>	27398,
		34486	=>	27395,
		34487	=>	27392,
		34488	=>	27388,
		34489	=>	27385,
		34490	=>	27382,
		34491	=>	27379,
		34492	=>	27376,
		34493	=>	27373,
		34494	=>	27370,
		34495	=>	27367,
		34496	=>	27364,
		34497	=>	27361,
		34498	=>	27358,
		34499	=>	27354,
		34500	=>	27351,
		34501	=>	27348,
		34502	=>	27345,
		34503	=>	27342,
		34504	=>	27339,
		34505	=>	27336,
		34506	=>	27333,
		34507	=>	27330,
		34508	=>	27327,
		34509	=>	27323,
		34510	=>	27320,
		34511	=>	27317,
		34512	=>	27314,
		34513	=>	27311,
		34514	=>	27308,
		34515	=>	27305,
		34516	=>	27302,
		34517	=>	27299,
		34518	=>	27296,
		34519	=>	27292,
		34520	=>	27289,
		34521	=>	27286,
		34522	=>	27283,
		34523	=>	27280,
		34524	=>	27277,
		34525	=>	27274,
		34526	=>	27271,
		34527	=>	27268,
		34528	=>	27265,
		34529	=>	27261,
		34530	=>	27258,
		34531	=>	27255,
		34532	=>	27252,
		34533	=>	27249,
		34534	=>	27246,
		34535	=>	27243,
		34536	=>	27240,
		34537	=>	27237,
		34538	=>	27234,
		34539	=>	27231,
		34540	=>	27227,
		34541	=>	27224,
		34542	=>	27221,
		34543	=>	27218,
		34544	=>	27215,
		34545	=>	27212,
		34546	=>	27209,
		34547	=>	27206,
		34548	=>	27203,
		34549	=>	27200,
		34550	=>	27196,
		34551	=>	27193,
		34552	=>	27190,
		34553	=>	27187,
		34554	=>	27184,
		34555	=>	27181,
		34556	=>	27178,
		34557	=>	27175,
		34558	=>	27172,
		34559	=>	27169,
		34560	=>	27166,
		34561	=>	27162,
		34562	=>	27159,
		34563	=>	27156,
		34564	=>	27153,
		34565	=>	27150,
		34566	=>	27147,
		34567	=>	27144,
		34568	=>	27141,
		34569	=>	27138,
		34570	=>	27135,
		34571	=>	27131,
		34572	=>	27128,
		34573	=>	27125,
		34574	=>	27122,
		34575	=>	27119,
		34576	=>	27116,
		34577	=>	27113,
		34578	=>	27110,
		34579	=>	27107,
		34580	=>	27104,
		34581	=>	27101,
		34582	=>	27097,
		34583	=>	27094,
		34584	=>	27091,
		34585	=>	27088,
		34586	=>	27085,
		34587	=>	27082,
		34588	=>	27079,
		34589	=>	27076,
		34590	=>	27073,
		34591	=>	27070,
		34592	=>	27066,
		34593	=>	27063,
		34594	=>	27060,
		34595	=>	27057,
		34596	=>	27054,
		34597	=>	27051,
		34598	=>	27048,
		34599	=>	27045,
		34600	=>	27042,
		34601	=>	27039,
		34602	=>	27036,
		34603	=>	27032,
		34604	=>	27029,
		34605	=>	27026,
		34606	=>	27023,
		34607	=>	27020,
		34608	=>	27017,
		34609	=>	27014,
		34610	=>	27011,
		34611	=>	27008,
		34612	=>	27005,
		34613	=>	27002,
		34614	=>	26998,
		34615	=>	26995,
		34616	=>	26992,
		34617	=>	26989,
		34618	=>	26986,
		34619	=>	26983,
		34620	=>	26980,
		34621	=>	26977,
		34622	=>	26974,
		34623	=>	26971,
		34624	=>	26968,
		34625	=>	26964,
		34626	=>	26961,
		34627	=>	26958,
		34628	=>	26955,
		34629	=>	26952,
		34630	=>	26949,
		34631	=>	26946,
		34632	=>	26943,
		34633	=>	26940,
		34634	=>	26937,
		34635	=>	26934,
		34636	=>	26930,
		34637	=>	26927,
		34638	=>	26924,
		34639	=>	26921,
		34640	=>	26918,
		34641	=>	26915,
		34642	=>	26912,
		34643	=>	26909,
		34644	=>	26906,
		34645	=>	26903,
		34646	=>	26900,
		34647	=>	26896,
		34648	=>	26893,
		34649	=>	26890,
		34650	=>	26887,
		34651	=>	26884,
		34652	=>	26881,
		34653	=>	26878,
		34654	=>	26875,
		34655	=>	26872,
		34656	=>	26869,
		34657	=>	26866,
		34658	=>	26862,
		34659	=>	26859,
		34660	=>	26856,
		34661	=>	26853,
		34662	=>	26850,
		34663	=>	26847,
		34664	=>	26844,
		34665	=>	26841,
		34666	=>	26838,
		34667	=>	26835,
		34668	=>	26832,
		34669	=>	26828,
		34670	=>	26825,
		34671	=>	26822,
		34672	=>	26819,
		34673	=>	26816,
		34674	=>	26813,
		34675	=>	26810,
		34676	=>	26807,
		34677	=>	26804,
		34678	=>	26801,
		34679	=>	26798,
		34680	=>	26794,
		34681	=>	26791,
		34682	=>	26788,
		34683	=>	26785,
		34684	=>	26782,
		34685	=>	26779,
		34686	=>	26776,
		34687	=>	26773,
		34688	=>	26770,
		34689	=>	26767,
		34690	=>	26764,
		34691	=>	26760,
		34692	=>	26757,
		34693	=>	26754,
		34694	=>	26751,
		34695	=>	26748,
		34696	=>	26745,
		34697	=>	26742,
		34698	=>	26739,
		34699	=>	26736,
		34700	=>	26733,
		34701	=>	26730,
		34702	=>	26727,
		34703	=>	26723,
		34704	=>	26720,
		34705	=>	26717,
		34706	=>	26714,
		34707	=>	26711,
		34708	=>	26708,
		34709	=>	26705,
		34710	=>	26702,
		34711	=>	26699,
		34712	=>	26696,
		34713	=>	26693,
		34714	=>	26689,
		34715	=>	26686,
		34716	=>	26683,
		34717	=>	26680,
		34718	=>	26677,
		34719	=>	26674,
		34720	=>	26671,
		34721	=>	26668,
		34722	=>	26665,
		34723	=>	26662,
		34724	=>	26659,
		34725	=>	26656,
		34726	=>	26652,
		34727	=>	26649,
		34728	=>	26646,
		34729	=>	26643,
		34730	=>	26640,
		34731	=>	26637,
		34732	=>	26634,
		34733	=>	26631,
		34734	=>	26628,
		34735	=>	26625,
		34736	=>	26622,
		34737	=>	26618,
		34738	=>	26615,
		34739	=>	26612,
		34740	=>	26609,
		34741	=>	26606,
		34742	=>	26603,
		34743	=>	26600,
		34744	=>	26597,
		34745	=>	26594,
		34746	=>	26591,
		34747	=>	26588,
		34748	=>	26585,
		34749	=>	26581,
		34750	=>	26578,
		34751	=>	26575,
		34752	=>	26572,
		34753	=>	26569,
		34754	=>	26566,
		34755	=>	26563,
		34756	=>	26560,
		34757	=>	26557,
		34758	=>	26554,
		34759	=>	26551,
		34760	=>	26548,
		34761	=>	26544,
		34762	=>	26541,
		34763	=>	26538,
		34764	=>	26535,
		34765	=>	26532,
		34766	=>	26529,
		34767	=>	26526,
		34768	=>	26523,
		34769	=>	26520,
		34770	=>	26517,
		34771	=>	26514,
		34772	=>	26511,
		34773	=>	26507,
		34774	=>	26504,
		34775	=>	26501,
		34776	=>	26498,
		34777	=>	26495,
		34778	=>	26492,
		34779	=>	26489,
		34780	=>	26486,
		34781	=>	26483,
		34782	=>	26480,
		34783	=>	26477,
		34784	=>	26474,
		34785	=>	26470,
		34786	=>	26467,
		34787	=>	26464,
		34788	=>	26461,
		34789	=>	26458,
		34790	=>	26455,
		34791	=>	26452,
		34792	=>	26449,
		34793	=>	26446,
		34794	=>	26443,
		34795	=>	26440,
		34796	=>	26437,
		34797	=>	26433,
		34798	=>	26430,
		34799	=>	26427,
		34800	=>	26424,
		34801	=>	26421,
		34802	=>	26418,
		34803	=>	26415,
		34804	=>	26412,
		34805	=>	26409,
		34806	=>	26406,
		34807	=>	26403,
		34808	=>	26400,
		34809	=>	26396,
		34810	=>	26393,
		34811	=>	26390,
		34812	=>	26387,
		34813	=>	26384,
		34814	=>	26381,
		34815	=>	26378,
		34816	=>	26375,
		34817	=>	26372,
		34818	=>	26369,
		34819	=>	26366,
		34820	=>	26363,
		34821	=>	26359,
		34822	=>	26356,
		34823	=>	26353,
		34824	=>	26350,
		34825	=>	26347,
		34826	=>	26344,
		34827	=>	26341,
		34828	=>	26338,
		34829	=>	26335,
		34830	=>	26332,
		34831	=>	26329,
		34832	=>	26326,
		34833	=>	26323,
		34834	=>	26319,
		34835	=>	26316,
		34836	=>	26313,
		34837	=>	26310,
		34838	=>	26307,
		34839	=>	26304,
		34840	=>	26301,
		34841	=>	26298,
		34842	=>	26295,
		34843	=>	26292,
		34844	=>	26289,
		34845	=>	26286,
		34846	=>	26282,
		34847	=>	26279,
		34848	=>	26276,
		34849	=>	26273,
		34850	=>	26270,
		34851	=>	26267,
		34852	=>	26264,
		34853	=>	26261,
		34854	=>	26258,
		34855	=>	26255,
		34856	=>	26252,
		34857	=>	26249,
		34858	=>	26246,
		34859	=>	26242,
		34860	=>	26239,
		34861	=>	26236,
		34862	=>	26233,
		34863	=>	26230,
		34864	=>	26227,
		34865	=>	26224,
		34866	=>	26221,
		34867	=>	26218,
		34868	=>	26215,
		34869	=>	26212,
		34870	=>	26209,
		34871	=>	26206,
		34872	=>	26202,
		34873	=>	26199,
		34874	=>	26196,
		34875	=>	26193,
		34876	=>	26190,
		34877	=>	26187,
		34878	=>	26184,
		34879	=>	26181,
		34880	=>	26178,
		34881	=>	26175,
		34882	=>	26172,
		34883	=>	26169,
		34884	=>	26165,
		34885	=>	26162,
		34886	=>	26159,
		34887	=>	26156,
		34888	=>	26153,
		34889	=>	26150,
		34890	=>	26147,
		34891	=>	26144,
		34892	=>	26141,
		34893	=>	26138,
		34894	=>	26135,
		34895	=>	26132,
		34896	=>	26129,
		34897	=>	26125,
		34898	=>	26122,
		34899	=>	26119,
		34900	=>	26116,
		34901	=>	26113,
		34902	=>	26110,
		34903	=>	26107,
		34904	=>	26104,
		34905	=>	26101,
		34906	=>	26098,
		34907	=>	26095,
		34908	=>	26092,
		34909	=>	26089,
		34910	=>	26086,
		34911	=>	26082,
		34912	=>	26079,
		34913	=>	26076,
		34914	=>	26073,
		34915	=>	26070,
		34916	=>	26067,
		34917	=>	26064,
		34918	=>	26061,
		34919	=>	26058,
		34920	=>	26055,
		34921	=>	26052,
		34922	=>	26049,
		34923	=>	26046,
		34924	=>	26042,
		34925	=>	26039,
		34926	=>	26036,
		34927	=>	26033,
		34928	=>	26030,
		34929	=>	26027,
		34930	=>	26024,
		34931	=>	26021,
		34932	=>	26018,
		34933	=>	26015,
		34934	=>	26012,
		34935	=>	26009,
		34936	=>	26006,
		34937	=>	26002,
		34938	=>	25999,
		34939	=>	25996,
		34940	=>	25993,
		34941	=>	25990,
		34942	=>	25987,
		34943	=>	25984,
		34944	=>	25981,
		34945	=>	25978,
		34946	=>	25975,
		34947	=>	25972,
		34948	=>	25969,
		34949	=>	25966,
		34950	=>	25963,
		34951	=>	25959,
		34952	=>	25956,
		34953	=>	25953,
		34954	=>	25950,
		34955	=>	25947,
		34956	=>	25944,
		34957	=>	25941,
		34958	=>	25938,
		34959	=>	25935,
		34960	=>	25932,
		34961	=>	25929,
		34962	=>	25926,
		34963	=>	25923,
		34964	=>	25920,
		34965	=>	25916,
		34966	=>	25913,
		34967	=>	25910,
		34968	=>	25907,
		34969	=>	25904,
		34970	=>	25901,
		34971	=>	25898,
		34972	=>	25895,
		34973	=>	25892,
		34974	=>	25889,
		34975	=>	25886,
		34976	=>	25883,
		34977	=>	25880,
		34978	=>	25877,
		34979	=>	25873,
		34980	=>	25870,
		34981	=>	25867,
		34982	=>	25864,
		34983	=>	25861,
		34984	=>	25858,
		34985	=>	25855,
		34986	=>	25852,
		34987	=>	25849,
		34988	=>	25846,
		34989	=>	25843,
		34990	=>	25840,
		34991	=>	25837,
		34992	=>	25834,
		34993	=>	25830,
		34994	=>	25827,
		34995	=>	25824,
		34996	=>	25821,
		34997	=>	25818,
		34998	=>	25815,
		34999	=>	25812,
		35000	=>	25809,
		35001	=>	25806,
		35002	=>	25803,
		35003	=>	25800,
		35004	=>	25797,
		35005	=>	25794,
		35006	=>	25791,
		35007	=>	25787,
		35008	=>	25784,
		35009	=>	25781,
		35010	=>	25778,
		35011	=>	25775,
		35012	=>	25772,
		35013	=>	25769,
		35014	=>	25766,
		35015	=>	25763,
		35016	=>	25760,
		35017	=>	25757,
		35018	=>	25754,
		35019	=>	25751,
		35020	=>	25748,
		35021	=>	25745,
		35022	=>	25741,
		35023	=>	25738,
		35024	=>	25735,
		35025	=>	25732,
		35026	=>	25729,
		35027	=>	25726,
		35028	=>	25723,
		35029	=>	25720,
		35030	=>	25717,
		35031	=>	25714,
		35032	=>	25711,
		35033	=>	25708,
		35034	=>	25705,
		35035	=>	25702,
		35036	=>	25698,
		35037	=>	25695,
		35038	=>	25692,
		35039	=>	25689,
		35040	=>	25686,
		35041	=>	25683,
		35042	=>	25680,
		35043	=>	25677,
		35044	=>	25674,
		35045	=>	25671,
		35046	=>	25668,
		35047	=>	25665,
		35048	=>	25662,
		35049	=>	25659,
		35050	=>	25656,
		35051	=>	25652,
		35052	=>	25649,
		35053	=>	25646,
		35054	=>	25643,
		35055	=>	25640,
		35056	=>	25637,
		35057	=>	25634,
		35058	=>	25631,
		35059	=>	25628,
		35060	=>	25625,
		35061	=>	25622,
		35062	=>	25619,
		35063	=>	25616,
		35064	=>	25613,
		35065	=>	25610,
		35066	=>	25606,
		35067	=>	25603,
		35068	=>	25600,
		35069	=>	25597,
		35070	=>	25594,
		35071	=>	25591,
		35072	=>	25588,
		35073	=>	25585,
		35074	=>	25582,
		35075	=>	25579,
		35076	=>	25576,
		35077	=>	25573,
		35078	=>	25570,
		35079	=>	25567,
		35080	=>	25564,
		35081	=>	25561,
		35082	=>	25557,
		35083	=>	25554,
		35084	=>	25551,
		35085	=>	25548,
		35086	=>	25545,
		35087	=>	25542,
		35088	=>	25539,
		35089	=>	25536,
		35090	=>	25533,
		35091	=>	25530,
		35092	=>	25527,
		35093	=>	25524,
		35094	=>	25521,
		35095	=>	25518,
		35096	=>	25515,
		35097	=>	25511,
		35098	=>	25508,
		35099	=>	25505,
		35100	=>	25502,
		35101	=>	25499,
		35102	=>	25496,
		35103	=>	25493,
		35104	=>	25490,
		35105	=>	25487,
		35106	=>	25484,
		35107	=>	25481,
		35108	=>	25478,
		35109	=>	25475,
		35110	=>	25472,
		35111	=>	25469,
		35112	=>	25466,
		35113	=>	25462,
		35114	=>	25459,
		35115	=>	25456,
		35116	=>	25453,
		35117	=>	25450,
		35118	=>	25447,
		35119	=>	25444,
		35120	=>	25441,
		35121	=>	25438,
		35122	=>	25435,
		35123	=>	25432,
		35124	=>	25429,
		35125	=>	25426,
		35126	=>	25423,
		35127	=>	25420,
		35128	=>	25417,
		35129	=>	25413,
		35130	=>	25410,
		35131	=>	25407,
		35132	=>	25404,
		35133	=>	25401,
		35134	=>	25398,
		35135	=>	25395,
		35136	=>	25392,
		35137	=>	25389,
		35138	=>	25386,
		35139	=>	25383,
		35140	=>	25380,
		35141	=>	25377,
		35142	=>	25374,
		35143	=>	25371,
		35144	=>	25368,
		35145	=>	25365,
		35146	=>	25361,
		35147	=>	25358,
		35148	=>	25355,
		35149	=>	25352,
		35150	=>	25349,
		35151	=>	25346,
		35152	=>	25343,
		35153	=>	25340,
		35154	=>	25337,
		35155	=>	25334,
		35156	=>	25331,
		35157	=>	25328,
		35158	=>	25325,
		35159	=>	25322,
		35160	=>	25319,
		35161	=>	25316,
		35162	=>	25313,
		35163	=>	25309,
		35164	=>	25306,
		35165	=>	25303,
		35166	=>	25300,
		35167	=>	25297,
		35168	=>	25294,
		35169	=>	25291,
		35170	=>	25288,
		35171	=>	25285,
		35172	=>	25282,
		35173	=>	25279,
		35174	=>	25276,
		35175	=>	25273,
		35176	=>	25270,
		35177	=>	25267,
		35178	=>	25264,
		35179	=>	25261,
		35180	=>	25257,
		35181	=>	25254,
		35182	=>	25251,
		35183	=>	25248,
		35184	=>	25245,
		35185	=>	25242,
		35186	=>	25239,
		35187	=>	25236,
		35188	=>	25233,
		35189	=>	25230,
		35190	=>	25227,
		35191	=>	25224,
		35192	=>	25221,
		35193	=>	25218,
		35194	=>	25215,
		35195	=>	25212,
		35196	=>	25209,
		35197	=>	25205,
		35198	=>	25202,
		35199	=>	25199,
		35200	=>	25196,
		35201	=>	25193,
		35202	=>	25190,
		35203	=>	25187,
		35204	=>	25184,
		35205	=>	25181,
		35206	=>	25178,
		35207	=>	25175,
		35208	=>	25172,
		35209	=>	25169,
		35210	=>	25166,
		35211	=>	25163,
		35212	=>	25160,
		35213	=>	25157,
		35214	=>	25154,
		35215	=>	25150,
		35216	=>	25147,
		35217	=>	25144,
		35218	=>	25141,
		35219	=>	25138,
		35220	=>	25135,
		35221	=>	25132,
		35222	=>	25129,
		35223	=>	25126,
		35224	=>	25123,
		35225	=>	25120,
		35226	=>	25117,
		35227	=>	25114,
		35228	=>	25111,
		35229	=>	25108,
		35230	=>	25105,
		35231	=>	25102,
		35232	=>	25099,
		35233	=>	25095,
		35234	=>	25092,
		35235	=>	25089,
		35236	=>	25086,
		35237	=>	25083,
		35238	=>	25080,
		35239	=>	25077,
		35240	=>	25074,
		35241	=>	25071,
		35242	=>	25068,
		35243	=>	25065,
		35244	=>	25062,
		35245	=>	25059,
		35246	=>	25056,
		35247	=>	25053,
		35248	=>	25050,
		35249	=>	25047,
		35250	=>	25044,
		35251	=>	25041,
		35252	=>	25037,
		35253	=>	25034,
		35254	=>	25031,
		35255	=>	25028,
		35256	=>	25025,
		35257	=>	25022,
		35258	=>	25019,
		35259	=>	25016,
		35260	=>	25013,
		35261	=>	25010,
		35262	=>	25007,
		35263	=>	25004,
		35264	=>	25001,
		35265	=>	24998,
		35266	=>	24995,
		35267	=>	24992,
		35268	=>	24989,
		35269	=>	24986,
		35270	=>	24983,
		35271	=>	24979,
		35272	=>	24976,
		35273	=>	24973,
		35274	=>	24970,
		35275	=>	24967,
		35276	=>	24964,
		35277	=>	24961,
		35278	=>	24958,
		35279	=>	24955,
		35280	=>	24952,
		35281	=>	24949,
		35282	=>	24946,
		35283	=>	24943,
		35284	=>	24940,
		35285	=>	24937,
		35286	=>	24934,
		35287	=>	24931,
		35288	=>	24928,
		35289	=>	24925,
		35290	=>	24922,
		35291	=>	24918,
		35292	=>	24915,
		35293	=>	24912,
		35294	=>	24909,
		35295	=>	24906,
		35296	=>	24903,
		35297	=>	24900,
		35298	=>	24897,
		35299	=>	24894,
		35300	=>	24891,
		35301	=>	24888,
		35302	=>	24885,
		35303	=>	24882,
		35304	=>	24879,
		35305	=>	24876,
		35306	=>	24873,
		35307	=>	24870,
		35308	=>	24867,
		35309	=>	24864,
		35310	=>	24861,
		35311	=>	24857,
		35312	=>	24854,
		35313	=>	24851,
		35314	=>	24848,
		35315	=>	24845,
		35316	=>	24842,
		35317	=>	24839,
		35318	=>	24836,
		35319	=>	24833,
		35320	=>	24830,
		35321	=>	24827,
		35322	=>	24824,
		35323	=>	24821,
		35324	=>	24818,
		35325	=>	24815,
		35326	=>	24812,
		35327	=>	24809,
		35328	=>	24806,
		35329	=>	24803,
		35330	=>	24800,
		35331	=>	24797,
		35332	=>	24793,
		35333	=>	24790,
		35334	=>	24787,
		35335	=>	24784,
		35336	=>	24781,
		35337	=>	24778,
		35338	=>	24775,
		35339	=>	24772,
		35340	=>	24769,
		35341	=>	24766,
		35342	=>	24763,
		35343	=>	24760,
		35344	=>	24757,
		35345	=>	24754,
		35346	=>	24751,
		35347	=>	24748,
		35348	=>	24745,
		35349	=>	24742,
		35350	=>	24739,
		35351	=>	24736,
		35352	=>	24733,
		35353	=>	24729,
		35354	=>	24726,
		35355	=>	24723,
		35356	=>	24720,
		35357	=>	24717,
		35358	=>	24714,
		35359	=>	24711,
		35360	=>	24708,
		35361	=>	24705,
		35362	=>	24702,
		35363	=>	24699,
		35364	=>	24696,
		35365	=>	24693,
		35366	=>	24690,
		35367	=>	24687,
		35368	=>	24684,
		35369	=>	24681,
		35370	=>	24678,
		35371	=>	24675,
		35372	=>	24672,
		35373	=>	24669,
		35374	=>	24666,
		35375	=>	24663,
		35376	=>	24659,
		35377	=>	24656,
		35378	=>	24653,
		35379	=>	24650,
		35380	=>	24647,
		35381	=>	24644,
		35382	=>	24641,
		35383	=>	24638,
		35384	=>	24635,
		35385	=>	24632,
		35386	=>	24629,
		35387	=>	24626,
		35388	=>	24623,
		35389	=>	24620,
		35390	=>	24617,
		35391	=>	24614,
		35392	=>	24611,
		35393	=>	24608,
		35394	=>	24605,
		35395	=>	24602,
		35396	=>	24599,
		35397	=>	24596,
		35398	=>	24593,
		35399	=>	24589,
		35400	=>	24586,
		35401	=>	24583,
		35402	=>	24580,
		35403	=>	24577,
		35404	=>	24574,
		35405	=>	24571,
		35406	=>	24568,
		35407	=>	24565,
		35408	=>	24562,
		35409	=>	24559,
		35410	=>	24556,
		35411	=>	24553,
		35412	=>	24550,
		35413	=>	24547,
		35414	=>	24544,
		35415	=>	24541,
		35416	=>	24538,
		35417	=>	24535,
		35418	=>	24532,
		35419	=>	24529,
		35420	=>	24526,
		35421	=>	24523,
		35422	=>	24520,
		35423	=>	24516,
		35424	=>	24513,
		35425	=>	24510,
		35426	=>	24507,
		35427	=>	24504,
		35428	=>	24501,
		35429	=>	24498,
		35430	=>	24495,
		35431	=>	24492,
		35432	=>	24489,
		35433	=>	24486,
		35434	=>	24483,
		35435	=>	24480,
		35436	=>	24477,
		35437	=>	24474,
		35438	=>	24471,
		35439	=>	24468,
		35440	=>	24465,
		35441	=>	24462,
		35442	=>	24459,
		35443	=>	24456,
		35444	=>	24453,
		35445	=>	24450,
		35446	=>	24447,
		35447	=>	24444,
		35448	=>	24440,
		35449	=>	24437,
		35450	=>	24434,
		35451	=>	24431,
		35452	=>	24428,
		35453	=>	24425,
		35454	=>	24422,
		35455	=>	24419,
		35456	=>	24416,
		35457	=>	24413,
		35458	=>	24410,
		35459	=>	24407,
		35460	=>	24404,
		35461	=>	24401,
		35462	=>	24398,
		35463	=>	24395,
		35464	=>	24392,
		35465	=>	24389,
		35466	=>	24386,
		35467	=>	24383,
		35468	=>	24380,
		35469	=>	24377,
		35470	=>	24374,
		35471	=>	24371,
		35472	=>	24368,
		35473	=>	24365,
		35474	=>	24362,
		35475	=>	24358,
		35476	=>	24355,
		35477	=>	24352,
		35478	=>	24349,
		35479	=>	24346,
		35480	=>	24343,
		35481	=>	24340,
		35482	=>	24337,
		35483	=>	24334,
		35484	=>	24331,
		35485	=>	24328,
		35486	=>	24325,
		35487	=>	24322,
		35488	=>	24319,
		35489	=>	24316,
		35490	=>	24313,
		35491	=>	24310,
		35492	=>	24307,
		35493	=>	24304,
		35494	=>	24301,
		35495	=>	24298,
		35496	=>	24295,
		35497	=>	24292,
		35498	=>	24289,
		35499	=>	24286,
		35500	=>	24283,
		35501	=>	24280,
		35502	=>	24277,
		35503	=>	24273,
		35504	=>	24270,
		35505	=>	24267,
		35506	=>	24264,
		35507	=>	24261,
		35508	=>	24258,
		35509	=>	24255,
		35510	=>	24252,
		35511	=>	24249,
		35512	=>	24246,
		35513	=>	24243,
		35514	=>	24240,
		35515	=>	24237,
		35516	=>	24234,
		35517	=>	24231,
		35518	=>	24228,
		35519	=>	24225,
		35520	=>	24222,
		35521	=>	24219,
		35522	=>	24216,
		35523	=>	24213,
		35524	=>	24210,
		35525	=>	24207,
		35526	=>	24204,
		35527	=>	24201,
		35528	=>	24198,
		35529	=>	24195,
		35530	=>	24192,
		35531	=>	24189,
		35532	=>	24186,
		35533	=>	24183,
		35534	=>	24179,
		35535	=>	24176,
		35536	=>	24173,
		35537	=>	24170,
		35538	=>	24167,
		35539	=>	24164,
		35540	=>	24161,
		35541	=>	24158,
		35542	=>	24155,
		35543	=>	24152,
		35544	=>	24149,
		35545	=>	24146,
		35546	=>	24143,
		35547	=>	24140,
		35548	=>	24137,
		35549	=>	24134,
		35550	=>	24131,
		35551	=>	24128,
		35552	=>	24125,
		35553	=>	24122,
		35554	=>	24119,
		35555	=>	24116,
		35556	=>	24113,
		35557	=>	24110,
		35558	=>	24107,
		35559	=>	24104,
		35560	=>	24101,
		35561	=>	24098,
		35562	=>	24095,
		35563	=>	24092,
		35564	=>	24089,
		35565	=>	24086,
		35566	=>	24083,
		35567	=>	24079,
		35568	=>	24076,
		35569	=>	24073,
		35570	=>	24070,
		35571	=>	24067,
		35572	=>	24064,
		35573	=>	24061,
		35574	=>	24058,
		35575	=>	24055,
		35576	=>	24052,
		35577	=>	24049,
		35578	=>	24046,
		35579	=>	24043,
		35580	=>	24040,
		35581	=>	24037,
		35582	=>	24034,
		35583	=>	24031,
		35584	=>	24028,
		35585	=>	24025,
		35586	=>	24022,
		35587	=>	24019,
		35588	=>	24016,
		35589	=>	24013,
		35590	=>	24010,
		35591	=>	24007,
		35592	=>	24004,
		35593	=>	24001,
		35594	=>	23998,
		35595	=>	23995,
		35596	=>	23992,
		35597	=>	23989,
		35598	=>	23986,
		35599	=>	23983,
		35600	=>	23980,
		35601	=>	23977,
		35602	=>	23974,
		35603	=>	23970,
		35604	=>	23967,
		35605	=>	23964,
		35606	=>	23961,
		35607	=>	23958,
		35608	=>	23955,
		35609	=>	23952,
		35610	=>	23949,
		35611	=>	23946,
		35612	=>	23943,
		35613	=>	23940,
		35614	=>	23937,
		35615	=>	23934,
		35616	=>	23931,
		35617	=>	23928,
		35618	=>	23925,
		35619	=>	23922,
		35620	=>	23919,
		35621	=>	23916,
		35622	=>	23913,
		35623	=>	23910,
		35624	=>	23907,
		35625	=>	23904,
		35626	=>	23901,
		35627	=>	23898,
		35628	=>	23895,
		35629	=>	23892,
		35630	=>	23889,
		35631	=>	23886,
		35632	=>	23883,
		35633	=>	23880,
		35634	=>	23877,
		35635	=>	23874,
		35636	=>	23871,
		35637	=>	23868,
		35638	=>	23865,
		35639	=>	23862,
		35640	=>	23859,
		35641	=>	23856,
		35642	=>	23853,
		35643	=>	23849,
		35644	=>	23846,
		35645	=>	23843,
		35646	=>	23840,
		35647	=>	23837,
		35648	=>	23834,
		35649	=>	23831,
		35650	=>	23828,
		35651	=>	23825,
		35652	=>	23822,
		35653	=>	23819,
		35654	=>	23816,
		35655	=>	23813,
		35656	=>	23810,
		35657	=>	23807,
		35658	=>	23804,
		35659	=>	23801,
		35660	=>	23798,
		35661	=>	23795,
		35662	=>	23792,
		35663	=>	23789,
		35664	=>	23786,
		35665	=>	23783,
		35666	=>	23780,
		35667	=>	23777,
		35668	=>	23774,
		35669	=>	23771,
		35670	=>	23768,
		35671	=>	23765,
		35672	=>	23762,
		35673	=>	23759,
		35674	=>	23756,
		35675	=>	23753,
		35676	=>	23750,
		35677	=>	23747,
		35678	=>	23744,
		35679	=>	23741,
		35680	=>	23738,
		35681	=>	23735,
		35682	=>	23732,
		35683	=>	23729,
		35684	=>	23726,
		35685	=>	23723,
		35686	=>	23720,
		35687	=>	23717,
		35688	=>	23714,
		35689	=>	23711,
		35690	=>	23708,
		35691	=>	23704,
		35692	=>	23701,
		35693	=>	23698,
		35694	=>	23695,
		35695	=>	23692,
		35696	=>	23689,
		35697	=>	23686,
		35698	=>	23683,
		35699	=>	23680,
		35700	=>	23677,
		35701	=>	23674,
		35702	=>	23671,
		35703	=>	23668,
		35704	=>	23665,
		35705	=>	23662,
		35706	=>	23659,
		35707	=>	23656,
		35708	=>	23653,
		35709	=>	23650,
		35710	=>	23647,
		35711	=>	23644,
		35712	=>	23641,
		35713	=>	23638,
		35714	=>	23635,
		35715	=>	23632,
		35716	=>	23629,
		35717	=>	23626,
		35718	=>	23623,
		35719	=>	23620,
		35720	=>	23617,
		35721	=>	23614,
		35722	=>	23611,
		35723	=>	23608,
		35724	=>	23605,
		35725	=>	23602,
		35726	=>	23599,
		35727	=>	23596,
		35728	=>	23593,
		35729	=>	23590,
		35730	=>	23587,
		35731	=>	23584,
		35732	=>	23581,
		35733	=>	23578,
		35734	=>	23575,
		35735	=>	23572,
		35736	=>	23569,
		35737	=>	23566,
		35738	=>	23563,
		35739	=>	23560,
		35740	=>	23557,
		35741	=>	23554,
		35742	=>	23551,
		35743	=>	23548,
		35744	=>	23545,
		35745	=>	23542,
		35746	=>	23539,
		35747	=>	23536,
		35748	=>	23533,
		35749	=>	23530,
		35750	=>	23527,
		35751	=>	23523,
		35752	=>	23520,
		35753	=>	23517,
		35754	=>	23514,
		35755	=>	23511,
		35756	=>	23508,
		35757	=>	23505,
		35758	=>	23502,
		35759	=>	23499,
		35760	=>	23496,
		35761	=>	23493,
		35762	=>	23490,
		35763	=>	23487,
		35764	=>	23484,
		35765	=>	23481,
		35766	=>	23478,
		35767	=>	23475,
		35768	=>	23472,
		35769	=>	23469,
		35770	=>	23466,
		35771	=>	23463,
		35772	=>	23460,
		35773	=>	23457,
		35774	=>	23454,
		35775	=>	23451,
		35776	=>	23448,
		35777	=>	23445,
		35778	=>	23442,
		35779	=>	23439,
		35780	=>	23436,
		35781	=>	23433,
		35782	=>	23430,
		35783	=>	23427,
		35784	=>	23424,
		35785	=>	23421,
		35786	=>	23418,
		35787	=>	23415,
		35788	=>	23412,
		35789	=>	23409,
		35790	=>	23406,
		35791	=>	23403,
		35792	=>	23400,
		35793	=>	23397,
		35794	=>	23394,
		35795	=>	23391,
		35796	=>	23388,
		35797	=>	23385,
		35798	=>	23382,
		35799	=>	23379,
		35800	=>	23376,
		35801	=>	23373,
		35802	=>	23370,
		35803	=>	23367,
		35804	=>	23364,
		35805	=>	23361,
		35806	=>	23358,
		35807	=>	23355,
		35808	=>	23352,
		35809	=>	23349,
		35810	=>	23346,
		35811	=>	23343,
		35812	=>	23340,
		35813	=>	23337,
		35814	=>	23334,
		35815	=>	23331,
		35816	=>	23328,
		35817	=>	23325,
		35818	=>	23322,
		35819	=>	23319,
		35820	=>	23316,
		35821	=>	23313,
		35822	=>	23310,
		35823	=>	23307,
		35824	=>	23304,
		35825	=>	23301,
		35826	=>	23298,
		35827	=>	23295,
		35828	=>	23292,
		35829	=>	23289,
		35830	=>	23286,
		35831	=>	23283,
		35832	=>	23280,
		35833	=>	23277,
		35834	=>	23274,
		35835	=>	23271,
		35836	=>	23268,
		35837	=>	23265,
		35838	=>	23262,
		35839	=>	23259,
		35840	=>	23256,
		35841	=>	23253,
		35842	=>	23250,
		35843	=>	23247,
		35844	=>	23244,
		35845	=>	23241,
		35846	=>	23238,
		35847	=>	23235,
		35848	=>	23232,
		35849	=>	23229,
		35850	=>	23226,
		35851	=>	23223,
		35852	=>	23220,
		35853	=>	23217,
		35854	=>	23214,
		35855	=>	23211,
		35856	=>	23208,
		35857	=>	23205,
		35858	=>	23201,
		35859	=>	23198,
		35860	=>	23195,
		35861	=>	23192,
		35862	=>	23189,
		35863	=>	23186,
		35864	=>	23183,
		35865	=>	23180,
		35866	=>	23177,
		35867	=>	23174,
		35868	=>	23171,
		35869	=>	23168,
		35870	=>	23165,
		35871	=>	23162,
		35872	=>	23159,
		35873	=>	23156,
		35874	=>	23153,
		35875	=>	23150,
		35876	=>	23147,
		35877	=>	23144,
		35878	=>	23141,
		35879	=>	23138,
		35880	=>	23135,
		35881	=>	23132,
		35882	=>	23129,
		35883	=>	23126,
		35884	=>	23123,
		35885	=>	23120,
		35886	=>	23117,
		35887	=>	23114,
		35888	=>	23111,
		35889	=>	23108,
		35890	=>	23105,
		35891	=>	23102,
		35892	=>	23099,
		35893	=>	23096,
		35894	=>	23093,
		35895	=>	23090,
		35896	=>	23087,
		35897	=>	23084,
		35898	=>	23081,
		35899	=>	23078,
		35900	=>	23075,
		35901	=>	23072,
		35902	=>	23069,
		35903	=>	23066,
		35904	=>	23063,
		35905	=>	23060,
		35906	=>	23057,
		35907	=>	23054,
		35908	=>	23051,
		35909	=>	23048,
		35910	=>	23045,
		35911	=>	23042,
		35912	=>	23039,
		35913	=>	23036,
		35914	=>	23033,
		35915	=>	23030,
		35916	=>	23027,
		35917	=>	23024,
		35918	=>	23021,
		35919	=>	23018,
		35920	=>	23015,
		35921	=>	23012,
		35922	=>	23009,
		35923	=>	23006,
		35924	=>	23003,
		35925	=>	23000,
		35926	=>	22997,
		35927	=>	22994,
		35928	=>	22991,
		35929	=>	22988,
		35930	=>	22985,
		35931	=>	22982,
		35932	=>	22979,
		35933	=>	22976,
		35934	=>	22973,
		35935	=>	22970,
		35936	=>	22967,
		35937	=>	22964,
		35938	=>	22961,
		35939	=>	22958,
		35940	=>	22955,
		35941	=>	22952,
		35942	=>	22949,
		35943	=>	22946,
		35944	=>	22943,
		35945	=>	22940,
		35946	=>	22937,
		35947	=>	22934,
		35948	=>	22931,
		35949	=>	22928,
		35950	=>	22925,
		35951	=>	22922,
		35952	=>	22919,
		35953	=>	22916,
		35954	=>	22913,
		35955	=>	22910,
		35956	=>	22907,
		35957	=>	22904,
		35958	=>	22901,
		35959	=>	22898,
		35960	=>	22895,
		35961	=>	22892,
		35962	=>	22889,
		35963	=>	22886,
		35964	=>	22884,
		35965	=>	22881,
		35966	=>	22878,
		35967	=>	22875,
		35968	=>	22872,
		35969	=>	22869,
		35970	=>	22866,
		35971	=>	22863,
		35972	=>	22860,
		35973	=>	22857,
		35974	=>	22854,
		35975	=>	22851,
		35976	=>	22848,
		35977	=>	22845,
		35978	=>	22842,
		35979	=>	22839,
		35980	=>	22836,
		35981	=>	22833,
		35982	=>	22830,
		35983	=>	22827,
		35984	=>	22824,
		35985	=>	22821,
		35986	=>	22818,
		35987	=>	22815,
		35988	=>	22812,
		35989	=>	22809,
		35990	=>	22806,
		35991	=>	22803,
		35992	=>	22800,
		35993	=>	22797,
		35994	=>	22794,
		35995	=>	22791,
		35996	=>	22788,
		35997	=>	22785,
		35998	=>	22782,
		35999	=>	22779,
		36000	=>	22776,
		36001	=>	22773,
		36002	=>	22770,
		36003	=>	22767,
		36004	=>	22764,
		36005	=>	22761,
		36006	=>	22758,
		36007	=>	22755,
		36008	=>	22752,
		36009	=>	22749,
		36010	=>	22746,
		36011	=>	22743,
		36012	=>	22740,
		36013	=>	22737,
		36014	=>	22734,
		36015	=>	22731,
		36016	=>	22728,
		36017	=>	22725,
		36018	=>	22722,
		36019	=>	22719,
		36020	=>	22716,
		36021	=>	22713,
		36022	=>	22710,
		36023	=>	22707,
		36024	=>	22704,
		36025	=>	22701,
		36026	=>	22698,
		36027	=>	22695,
		36028	=>	22692,
		36029	=>	22689,
		36030	=>	22686,
		36031	=>	22683,
		36032	=>	22680,
		36033	=>	22677,
		36034	=>	22674,
		36035	=>	22671,
		36036	=>	22668,
		36037	=>	22665,
		36038	=>	22662,
		36039	=>	22659,
		36040	=>	22656,
		36041	=>	22653,
		36042	=>	22650,
		36043	=>	22647,
		36044	=>	22644,
		36045	=>	22641,
		36046	=>	22638,
		36047	=>	22635,
		36048	=>	22632,
		36049	=>	22629,
		36050	=>	22626,
		36051	=>	22623,
		36052	=>	22620,
		36053	=>	22617,
		36054	=>	22614,
		36055	=>	22611,
		36056	=>	22608,
		36057	=>	22605,
		36058	=>	22602,
		36059	=>	22599,
		36060	=>	22596,
		36061	=>	22593,
		36062	=>	22590,
		36063	=>	22587,
		36064	=>	22584,
		36065	=>	22581,
		36066	=>	22578,
		36067	=>	22575,
		36068	=>	22572,
		36069	=>	22570,
		36070	=>	22567,
		36071	=>	22564,
		36072	=>	22561,
		36073	=>	22558,
		36074	=>	22555,
		36075	=>	22552,
		36076	=>	22549,
		36077	=>	22546,
		36078	=>	22543,
		36079	=>	22540,
		36080	=>	22537,
		36081	=>	22534,
		36082	=>	22531,
		36083	=>	22528,
		36084	=>	22525,
		36085	=>	22522,
		36086	=>	22519,
		36087	=>	22516,
		36088	=>	22513,
		36089	=>	22510,
		36090	=>	22507,
		36091	=>	22504,
		36092	=>	22501,
		36093	=>	22498,
		36094	=>	22495,
		36095	=>	22492,
		36096	=>	22489,
		36097	=>	22486,
		36098	=>	22483,
		36099	=>	22480,
		36100	=>	22477,
		36101	=>	22474,
		36102	=>	22471,
		36103	=>	22468,
		36104	=>	22465,
		36105	=>	22462,
		36106	=>	22459,
		36107	=>	22456,
		36108	=>	22453,
		36109	=>	22450,
		36110	=>	22447,
		36111	=>	22444,
		36112	=>	22441,
		36113	=>	22438,
		36114	=>	22435,
		36115	=>	22432,
		36116	=>	22429,
		36117	=>	22426,
		36118	=>	22423,
		36119	=>	22420,
		36120	=>	22417,
		36121	=>	22414,
		36122	=>	22411,
		36123	=>	22408,
		36124	=>	22405,
		36125	=>	22402,
		36126	=>	22399,
		36127	=>	22397,
		36128	=>	22394,
		36129	=>	22391,
		36130	=>	22388,
		36131	=>	22385,
		36132	=>	22382,
		36133	=>	22379,
		36134	=>	22376,
		36135	=>	22373,
		36136	=>	22370,
		36137	=>	22367,
		36138	=>	22364,
		36139	=>	22361,
		36140	=>	22358,
		36141	=>	22355,
		36142	=>	22352,
		36143	=>	22349,
		36144	=>	22346,
		36145	=>	22343,
		36146	=>	22340,
		36147	=>	22337,
		36148	=>	22334,
		36149	=>	22331,
		36150	=>	22328,
		36151	=>	22325,
		36152	=>	22322,
		36153	=>	22319,
		36154	=>	22316,
		36155	=>	22313,
		36156	=>	22310,
		36157	=>	22307,
		36158	=>	22304,
		36159	=>	22301,
		36160	=>	22298,
		36161	=>	22295,
		36162	=>	22292,
		36163	=>	22289,
		36164	=>	22286,
		36165	=>	22283,
		36166	=>	22280,
		36167	=>	22277,
		36168	=>	22274,
		36169	=>	22271,
		36170	=>	22268,
		36171	=>	22265,
		36172	=>	22263,
		36173	=>	22260,
		36174	=>	22257,
		36175	=>	22254,
		36176	=>	22251,
		36177	=>	22248,
		36178	=>	22245,
		36179	=>	22242,
		36180	=>	22239,
		36181	=>	22236,
		36182	=>	22233,
		36183	=>	22230,
		36184	=>	22227,
		36185	=>	22224,
		36186	=>	22221,
		36187	=>	22218,
		36188	=>	22215,
		36189	=>	22212,
		36190	=>	22209,
		36191	=>	22206,
		36192	=>	22203,
		36193	=>	22200,
		36194	=>	22197,
		36195	=>	22194,
		36196	=>	22191,
		36197	=>	22188,
		36198	=>	22185,
		36199	=>	22182,
		36200	=>	22179,
		36201	=>	22176,
		36202	=>	22173,
		36203	=>	22170,
		36204	=>	22167,
		36205	=>	22164,
		36206	=>	22161,
		36207	=>	22158,
		36208	=>	22155,
		36209	=>	22152,
		36210	=>	22149,
		36211	=>	22147,
		36212	=>	22144,
		36213	=>	22141,
		36214	=>	22138,
		36215	=>	22135,
		36216	=>	22132,
		36217	=>	22129,
		36218	=>	22126,
		36219	=>	22123,
		36220	=>	22120,
		36221	=>	22117,
		36222	=>	22114,
		36223	=>	22111,
		36224	=>	22108,
		36225	=>	22105,
		36226	=>	22102,
		36227	=>	22099,
		36228	=>	22096,
		36229	=>	22093,
		36230	=>	22090,
		36231	=>	22087,
		36232	=>	22084,
		36233	=>	22081,
		36234	=>	22078,
		36235	=>	22075,
		36236	=>	22072,
		36237	=>	22069,
		36238	=>	22066,
		36239	=>	22063,
		36240	=>	22060,
		36241	=>	22057,
		36242	=>	22054,
		36243	=>	22051,
		36244	=>	22049,
		36245	=>	22046,
		36246	=>	22043,
		36247	=>	22040,
		36248	=>	22037,
		36249	=>	22034,
		36250	=>	22031,
		36251	=>	22028,
		36252	=>	22025,
		36253	=>	22022,
		36254	=>	22019,
		36255	=>	22016,
		36256	=>	22013,
		36257	=>	22010,
		36258	=>	22007,
		36259	=>	22004,
		36260	=>	22001,
		36261	=>	21998,
		36262	=>	21995,
		36263	=>	21992,
		36264	=>	21989,
		36265	=>	21986,
		36266	=>	21983,
		36267	=>	21980,
		36268	=>	21977,
		36269	=>	21974,
		36270	=>	21971,
		36271	=>	21968,
		36272	=>	21965,
		36273	=>	21962,
		36274	=>	21959,
		36275	=>	21957,
		36276	=>	21954,
		36277	=>	21951,
		36278	=>	21948,
		36279	=>	21945,
		36280	=>	21942,
		36281	=>	21939,
		36282	=>	21936,
		36283	=>	21933,
		36284	=>	21930,
		36285	=>	21927,
		36286	=>	21924,
		36287	=>	21921,
		36288	=>	21918,
		36289	=>	21915,
		36290	=>	21912,
		36291	=>	21909,
		36292	=>	21906,
		36293	=>	21903,
		36294	=>	21900,
		36295	=>	21897,
		36296	=>	21894,
		36297	=>	21891,
		36298	=>	21888,
		36299	=>	21885,
		36300	=>	21882,
		36301	=>	21879,
		36302	=>	21876,
		36303	=>	21874,
		36304	=>	21871,
		36305	=>	21868,
		36306	=>	21865,
		36307	=>	21862,
		36308	=>	21859,
		36309	=>	21856,
		36310	=>	21853,
		36311	=>	21850,
		36312	=>	21847,
		36313	=>	21844,
		36314	=>	21841,
		36315	=>	21838,
		36316	=>	21835,
		36317	=>	21832,
		36318	=>	21829,
		36319	=>	21826,
		36320	=>	21823,
		36321	=>	21820,
		36322	=>	21817,
		36323	=>	21814,
		36324	=>	21811,
		36325	=>	21808,
		36326	=>	21805,
		36327	=>	21802,
		36328	=>	21799,
		36329	=>	21797,
		36330	=>	21794,
		36331	=>	21791,
		36332	=>	21788,
		36333	=>	21785,
		36334	=>	21782,
		36335	=>	21779,
		36336	=>	21776,
		36337	=>	21773,
		36338	=>	21770,
		36339	=>	21767,
		36340	=>	21764,
		36341	=>	21761,
		36342	=>	21758,
		36343	=>	21755,
		36344	=>	21752,
		36345	=>	21749,
		36346	=>	21746,
		36347	=>	21743,
		36348	=>	21740,
		36349	=>	21737,
		36350	=>	21734,
		36351	=>	21731,
		36352	=>	21728,
		36353	=>	21726,
		36354	=>	21723,
		36355	=>	21720,
		36356	=>	21717,
		36357	=>	21714,
		36358	=>	21711,
		36359	=>	21708,
		36360	=>	21705,
		36361	=>	21702,
		36362	=>	21699,
		36363	=>	21696,
		36364	=>	21693,
		36365	=>	21690,
		36366	=>	21687,
		36367	=>	21684,
		36368	=>	21681,
		36369	=>	21678,
		36370	=>	21675,
		36371	=>	21672,
		36372	=>	21669,
		36373	=>	21666,
		36374	=>	21663,
		36375	=>	21660,
		36376	=>	21658,
		36377	=>	21655,
		36378	=>	21652,
		36379	=>	21649,
		36380	=>	21646,
		36381	=>	21643,
		36382	=>	21640,
		36383	=>	21637,
		36384	=>	21634,
		36385	=>	21631,
		36386	=>	21628,
		36387	=>	21625,
		36388	=>	21622,
		36389	=>	21619,
		36390	=>	21616,
		36391	=>	21613,
		36392	=>	21610,
		36393	=>	21607,
		36394	=>	21604,
		36395	=>	21601,
		36396	=>	21598,
		36397	=>	21595,
		36398	=>	21593,
		36399	=>	21590,
		36400	=>	21587,
		36401	=>	21584,
		36402	=>	21581,
		36403	=>	21578,
		36404	=>	21575,
		36405	=>	21572,
		36406	=>	21569,
		36407	=>	21566,
		36408	=>	21563,
		36409	=>	21560,
		36410	=>	21557,
		36411	=>	21554,
		36412	=>	21551,
		36413	=>	21548,
		36414	=>	21545,
		36415	=>	21542,
		36416	=>	21539,
		36417	=>	21536,
		36418	=>	21533,
		36419	=>	21531,
		36420	=>	21528,
		36421	=>	21525,
		36422	=>	21522,
		36423	=>	21519,
		36424	=>	21516,
		36425	=>	21513,
		36426	=>	21510,
		36427	=>	21507,
		36428	=>	21504,
		36429	=>	21501,
		36430	=>	21498,
		36431	=>	21495,
		36432	=>	21492,
		36433	=>	21489,
		36434	=>	21486,
		36435	=>	21483,
		36436	=>	21480,
		36437	=>	21477,
		36438	=>	21474,
		36439	=>	21472,
		36440	=>	21469,
		36441	=>	21466,
		36442	=>	21463,
		36443	=>	21460,
		36444	=>	21457,
		36445	=>	21454,
		36446	=>	21451,
		36447	=>	21448,
		36448	=>	21445,
		36449	=>	21442,
		36450	=>	21439,
		36451	=>	21436,
		36452	=>	21433,
		36453	=>	21430,
		36454	=>	21427,
		36455	=>	21424,
		36456	=>	21421,
		36457	=>	21418,
		36458	=>	21415,
		36459	=>	21413,
		36460	=>	21410,
		36461	=>	21407,
		36462	=>	21404,
		36463	=>	21401,
		36464	=>	21398,
		36465	=>	21395,
		36466	=>	21392,
		36467	=>	21389,
		36468	=>	21386,
		36469	=>	21383,
		36470	=>	21380,
		36471	=>	21377,
		36472	=>	21374,
		36473	=>	21371,
		36474	=>	21368,
		36475	=>	21365,
		36476	=>	21362,
		36477	=>	21360,
		36478	=>	21357,
		36479	=>	21354,
		36480	=>	21351,
		36481	=>	21348,
		36482	=>	21345,
		36483	=>	21342,
		36484	=>	21339,
		36485	=>	21336,
		36486	=>	21333,
		36487	=>	21330,
		36488	=>	21327,
		36489	=>	21324,
		36490	=>	21321,
		36491	=>	21318,
		36492	=>	21315,
		36493	=>	21312,
		36494	=>	21309,
		36495	=>	21307,
		36496	=>	21304,
		36497	=>	21301,
		36498	=>	21298,
		36499	=>	21295,
		36500	=>	21292,
		36501	=>	21289,
		36502	=>	21286,
		36503	=>	21283,
		36504	=>	21280,
		36505	=>	21277,
		36506	=>	21274,
		36507	=>	21271,
		36508	=>	21268,
		36509	=>	21265,
		36510	=>	21262,
		36511	=>	21259,
		36512	=>	21257,
		36513	=>	21254,
		36514	=>	21251,
		36515	=>	21248,
		36516	=>	21245,
		36517	=>	21242,
		36518	=>	21239,
		36519	=>	21236,
		36520	=>	21233,
		36521	=>	21230,
		36522	=>	21227,
		36523	=>	21224,
		36524	=>	21221,
		36525	=>	21218,
		36526	=>	21215,
		36527	=>	21212,
		36528	=>	21209,
		36529	=>	21207,
		36530	=>	21204,
		36531	=>	21201,
		36532	=>	21198,
		36533	=>	21195,
		36534	=>	21192,
		36535	=>	21189,
		36536	=>	21186,
		36537	=>	21183,
		36538	=>	21180,
		36539	=>	21177,
		36540	=>	21174,
		36541	=>	21171,
		36542	=>	21168,
		36543	=>	21165,
		36544	=>	21162,
		36545	=>	21160,
		36546	=>	21157,
		36547	=>	21154,
		36548	=>	21151,
		36549	=>	21148,
		36550	=>	21145,
		36551	=>	21142,
		36552	=>	21139,
		36553	=>	21136,
		36554	=>	21133,
		36555	=>	21130,
		36556	=>	21127,
		36557	=>	21124,
		36558	=>	21121,
		36559	=>	21118,
		36560	=>	21115,
		36561	=>	21113,
		36562	=>	21110,
		36563	=>	21107,
		36564	=>	21104,
		36565	=>	21101,
		36566	=>	21098,
		36567	=>	21095,
		36568	=>	21092,
		36569	=>	21089,
		36570	=>	21086,
		36571	=>	21083,
		36572	=>	21080,
		36573	=>	21077,
		36574	=>	21074,
		36575	=>	21071,
		36576	=>	21068,
		36577	=>	21066,
		36578	=>	21063,
		36579	=>	21060,
		36580	=>	21057,
		36581	=>	21054,
		36582	=>	21051,
		36583	=>	21048,
		36584	=>	21045,
		36585	=>	21042,
		36586	=>	21039,
		36587	=>	21036,
		36588	=>	21033,
		36589	=>	21030,
		36590	=>	21027,
		36591	=>	21024,
		36592	=>	21022,
		36593	=>	21019,
		36594	=>	21016,
		36595	=>	21013,
		36596	=>	21010,
		36597	=>	21007,
		36598	=>	21004,
		36599	=>	21001,
		36600	=>	20998,
		36601	=>	20995,
		36602	=>	20992,
		36603	=>	20989,
		36604	=>	20986,
		36605	=>	20983,
		36606	=>	20981,
		36607	=>	20978,
		36608	=>	20975,
		36609	=>	20972,
		36610	=>	20969,
		36611	=>	20966,
		36612	=>	20963,
		36613	=>	20960,
		36614	=>	20957,
		36615	=>	20954,
		36616	=>	20951,
		36617	=>	20948,
		36618	=>	20945,
		36619	=>	20942,
		36620	=>	20939,
		36621	=>	20937,
		36622	=>	20934,
		36623	=>	20931,
		36624	=>	20928,
		36625	=>	20925,
		36626	=>	20922,
		36627	=>	20919,
		36628	=>	20916,
		36629	=>	20913,
		36630	=>	20910,
		36631	=>	20907,
		36632	=>	20904,
		36633	=>	20901,
		36634	=>	20898,
		36635	=>	20896,
		36636	=>	20893,
		36637	=>	20890,
		36638	=>	20887,
		36639	=>	20884,
		36640	=>	20881,
		36641	=>	20878,
		36642	=>	20875,
		36643	=>	20872,
		36644	=>	20869,
		36645	=>	20866,
		36646	=>	20863,
		36647	=>	20860,
		36648	=>	20857,
		36649	=>	20855,
		36650	=>	20852,
		36651	=>	20849,
		36652	=>	20846,
		36653	=>	20843,
		36654	=>	20840,
		36655	=>	20837,
		36656	=>	20834,
		36657	=>	20831,
		36658	=>	20828,
		36659	=>	20825,
		36660	=>	20822,
		36661	=>	20819,
		36662	=>	20817,
		36663	=>	20814,
		36664	=>	20811,
		36665	=>	20808,
		36666	=>	20805,
		36667	=>	20802,
		36668	=>	20799,
		36669	=>	20796,
		36670	=>	20793,
		36671	=>	20790,
		36672	=>	20787,
		36673	=>	20784,
		36674	=>	20781,
		36675	=>	20779,
		36676	=>	20776,
		36677	=>	20773,
		36678	=>	20770,
		36679	=>	20767,
		36680	=>	20764,
		36681	=>	20761,
		36682	=>	20758,
		36683	=>	20755,
		36684	=>	20752,
		36685	=>	20749,
		36686	=>	20746,
		36687	=>	20743,
		36688	=>	20741,
		36689	=>	20738,
		36690	=>	20735,
		36691	=>	20732,
		36692	=>	20729,
		36693	=>	20726,
		36694	=>	20723,
		36695	=>	20720,
		36696	=>	20717,
		36697	=>	20714,
		36698	=>	20711,
		36699	=>	20708,
		36700	=>	20705,
		36701	=>	20703,
		36702	=>	20700,
		36703	=>	20697,
		36704	=>	20694,
		36705	=>	20691,
		36706	=>	20688,
		36707	=>	20685,
		36708	=>	20682,
		36709	=>	20679,
		36710	=>	20676,
		36711	=>	20673,
		36712	=>	20670,
		36713	=>	20667,
		36714	=>	20665,
		36715	=>	20662,
		36716	=>	20659,
		36717	=>	20656,
		36718	=>	20653,
		36719	=>	20650,
		36720	=>	20647,
		36721	=>	20644,
		36722	=>	20641,
		36723	=>	20638,
		36724	=>	20635,
		36725	=>	20632,
		36726	=>	20630,
		36727	=>	20627,
		36728	=>	20624,
		36729	=>	20621,
		36730	=>	20618,
		36731	=>	20615,
		36732	=>	20612,
		36733	=>	20609,
		36734	=>	20606,
		36735	=>	20603,
		36736	=>	20600,
		36737	=>	20597,
		36738	=>	20595,
		36739	=>	20592,
		36740	=>	20589,
		36741	=>	20586,
		36742	=>	20583,
		36743	=>	20580,
		36744	=>	20577,
		36745	=>	20574,
		36746	=>	20571,
		36747	=>	20568,
		36748	=>	20565,
		36749	=>	20562,
		36750	=>	20560,
		36751	=>	20557,
		36752	=>	20554,
		36753	=>	20551,
		36754	=>	20548,
		36755	=>	20545,
		36756	=>	20542,
		36757	=>	20539,
		36758	=>	20536,
		36759	=>	20533,
		36760	=>	20530,
		36761	=>	20527,
		36762	=>	20525,
		36763	=>	20522,
		36764	=>	20519,
		36765	=>	20516,
		36766	=>	20513,
		36767	=>	20510,
		36768	=>	20507,
		36769	=>	20504,
		36770	=>	20501,
		36771	=>	20498,
		36772	=>	20495,
		36773	=>	20493,
		36774	=>	20490,
		36775	=>	20487,
		36776	=>	20484,
		36777	=>	20481,
		36778	=>	20478,
		36779	=>	20475,
		36780	=>	20472,
		36781	=>	20469,
		36782	=>	20466,
		36783	=>	20463,
		36784	=>	20460,
		36785	=>	20458,
		36786	=>	20455,
		36787	=>	20452,
		36788	=>	20449,
		36789	=>	20446,
		36790	=>	20443,
		36791	=>	20440,
		36792	=>	20437,
		36793	=>	20434,
		36794	=>	20431,
		36795	=>	20428,
		36796	=>	20426,
		36797	=>	20423,
		36798	=>	20420,
		36799	=>	20417,
		36800	=>	20414,
		36801	=>	20411,
		36802	=>	20408,
		36803	=>	20405,
		36804	=>	20402,
		36805	=>	20399,
		36806	=>	20396,
		36807	=>	20394,
		36808	=>	20391,
		36809	=>	20388,
		36810	=>	20385,
		36811	=>	20382,
		36812	=>	20379,
		36813	=>	20376,
		36814	=>	20373,
		36815	=>	20370,
		36816	=>	20367,
		36817	=>	20364,
		36818	=>	20362,
		36819	=>	20359,
		36820	=>	20356,
		36821	=>	20353,
		36822	=>	20350,
		36823	=>	20347,
		36824	=>	20344,
		36825	=>	20341,
		36826	=>	20338,
		36827	=>	20335,
		36828	=>	20332,
		36829	=>	20330,
		36830	=>	20327,
		36831	=>	20324,
		36832	=>	20321,
		36833	=>	20318,
		36834	=>	20315,
		36835	=>	20312,
		36836	=>	20309,
		36837	=>	20306,
		36838	=>	20303,
		36839	=>	20301,
		36840	=>	20298,
		36841	=>	20295,
		36842	=>	20292,
		36843	=>	20289,
		36844	=>	20286,
		36845	=>	20283,
		36846	=>	20280,
		36847	=>	20277,
		36848	=>	20274,
		36849	=>	20271,
		36850	=>	20269,
		36851	=>	20266,
		36852	=>	20263,
		36853	=>	20260,
		36854	=>	20257,
		36855	=>	20254,
		36856	=>	20251,
		36857	=>	20248,
		36858	=>	20245,
		36859	=>	20242,
		36860	=>	20240,
		36861	=>	20237,
		36862	=>	20234,
		36863	=>	20231,
		36864	=>	20228,
		36865	=>	20225,
		36866	=>	20222,
		36867	=>	20219,
		36868	=>	20216,
		36869	=>	20213,
		36870	=>	20211,
		36871	=>	20208,
		36872	=>	20205,
		36873	=>	20202,
		36874	=>	20199,
		36875	=>	20196,
		36876	=>	20193,
		36877	=>	20190,
		36878	=>	20187,
		36879	=>	20184,
		36880	=>	20181,
		36881	=>	20179,
		36882	=>	20176,
		36883	=>	20173,
		36884	=>	20170,
		36885	=>	20167,
		36886	=>	20164,
		36887	=>	20161,
		36888	=>	20158,
		36889	=>	20155,
		36890	=>	20152,
		36891	=>	20150,
		36892	=>	20147,
		36893	=>	20144,
		36894	=>	20141,
		36895	=>	20138,
		36896	=>	20135,
		36897	=>	20132,
		36898	=>	20129,
		36899	=>	20126,
		36900	=>	20124,
		36901	=>	20121,
		36902	=>	20118,
		36903	=>	20115,
		36904	=>	20112,
		36905	=>	20109,
		36906	=>	20106,
		36907	=>	20103,
		36908	=>	20100,
		36909	=>	20097,
		36910	=>	20095,
		36911	=>	20092,
		36912	=>	20089,
		36913	=>	20086,
		36914	=>	20083,
		36915	=>	20080,
		36916	=>	20077,
		36917	=>	20074,
		36918	=>	20071,
		36919	=>	20068,
		36920	=>	20066,
		36921	=>	20063,
		36922	=>	20060,
		36923	=>	20057,
		36924	=>	20054,
		36925	=>	20051,
		36926	=>	20048,
		36927	=>	20045,
		36928	=>	20042,
		36929	=>	20040,
		36930	=>	20037,
		36931	=>	20034,
		36932	=>	20031,
		36933	=>	20028,
		36934	=>	20025,
		36935	=>	20022,
		36936	=>	20019,
		36937	=>	20016,
		36938	=>	20013,
		36939	=>	20011,
		36940	=>	20008,
		36941	=>	20005,
		36942	=>	20002,
		36943	=>	19999,
		36944	=>	19996,
		36945	=>	19993,
		36946	=>	19990,
		36947	=>	19987,
		36948	=>	19985,
		36949	=>	19982,
		36950	=>	19979,
		36951	=>	19976,
		36952	=>	19973,
		36953	=>	19970,
		36954	=>	19967,
		36955	=>	19964,
		36956	=>	19961,
		36957	=>	19958,
		36958	=>	19956,
		36959	=>	19953,
		36960	=>	19950,
		36961	=>	19947,
		36962	=>	19944,
		36963	=>	19941,
		36964	=>	19938,
		36965	=>	19935,
		36966	=>	19932,
		36967	=>	19930,
		36968	=>	19927,
		36969	=>	19924,
		36970	=>	19921,
		36971	=>	19918,
		36972	=>	19915,
		36973	=>	19912,
		36974	=>	19909,
		36975	=>	19906,
		36976	=>	19904,
		36977	=>	19901,
		36978	=>	19898,
		36979	=>	19895,
		36980	=>	19892,
		36981	=>	19889,
		36982	=>	19886,
		36983	=>	19883,
		36984	=>	19880,
		36985	=>	19878,
		36986	=>	19875,
		36987	=>	19872,
		36988	=>	19869,
		36989	=>	19866,
		36990	=>	19863,
		36991	=>	19860,
		36992	=>	19857,
		36993	=>	19854,
		36994	=>	19852,
		36995	=>	19849,
		36996	=>	19846,
		36997	=>	19843,
		36998	=>	19840,
		36999	=>	19837,
		37000	=>	19834,
		37001	=>	19831,
		37002	=>	19828,
		37003	=>	19826,
		37004	=>	19823,
		37005	=>	19820,
		37006	=>	19817,
		37007	=>	19814,
		37008	=>	19811,
		37009	=>	19808,
		37010	=>	19805,
		37011	=>	19803,
		37012	=>	19800,
		37013	=>	19797,
		37014	=>	19794,
		37015	=>	19791,
		37016	=>	19788,
		37017	=>	19785,
		37018	=>	19782,
		37019	=>	19779,
		37020	=>	19777,
		37021	=>	19774,
		37022	=>	19771,
		37023	=>	19768,
		37024	=>	19765,
		37025	=>	19762,
		37026	=>	19759,
		37027	=>	19756,
		37028	=>	19753,
		37029	=>	19751,
		37030	=>	19748,
		37031	=>	19745,
		37032	=>	19742,
		37033	=>	19739,
		37034	=>	19736,
		37035	=>	19733,
		37036	=>	19730,
		37037	=>	19728,
		37038	=>	19725,
		37039	=>	19722,
		37040	=>	19719,
		37041	=>	19716,
		37042	=>	19713,
		37043	=>	19710,
		37044	=>	19707,
		37045	=>	19704,
		37046	=>	19702,
		37047	=>	19699,
		37048	=>	19696,
		37049	=>	19693,
		37050	=>	19690,
		37051	=>	19687,
		37052	=>	19684,
		37053	=>	19681,
		37054	=>	19679,
		37055	=>	19676,
		37056	=>	19673,
		37057	=>	19670,
		37058	=>	19667,
		37059	=>	19664,
		37060	=>	19661,
		37061	=>	19658,
		37062	=>	19656,
		37063	=>	19653,
		37064	=>	19650,
		37065	=>	19647,
		37066	=>	19644,
		37067	=>	19641,
		37068	=>	19638,
		37069	=>	19635,
		37070	=>	19633,
		37071	=>	19630,
		37072	=>	19627,
		37073	=>	19624,
		37074	=>	19621,
		37075	=>	19618,
		37076	=>	19615,
		37077	=>	19612,
		37078	=>	19609,
		37079	=>	19607,
		37080	=>	19604,
		37081	=>	19601,
		37082	=>	19598,
		37083	=>	19595,
		37084	=>	19592,
		37085	=>	19589,
		37086	=>	19586,
		37087	=>	19584,
		37088	=>	19581,
		37089	=>	19578,
		37090	=>	19575,
		37091	=>	19572,
		37092	=>	19569,
		37093	=>	19566,
		37094	=>	19563,
		37095	=>	19561,
		37096	=>	19558,
		37097	=>	19555,
		37098	=>	19552,
		37099	=>	19549,
		37100	=>	19546,
		37101	=>	19543,
		37102	=>	19540,
		37103	=>	19538,
		37104	=>	19535,
		37105	=>	19532,
		37106	=>	19529,
		37107	=>	19526,
		37108	=>	19523,
		37109	=>	19520,
		37110	=>	19517,
		37111	=>	19515,
		37112	=>	19512,
		37113	=>	19509,
		37114	=>	19506,
		37115	=>	19503,
		37116	=>	19500,
		37117	=>	19497,
		37118	=>	19494,
		37119	=>	19492,
		37120	=>	19489,
		37121	=>	19486,
		37122	=>	19483,
		37123	=>	19480,
		37124	=>	19477,
		37125	=>	19474,
		37126	=>	19472,
		37127	=>	19469,
		37128	=>	19466,
		37129	=>	19463,
		37130	=>	19460,
		37131	=>	19457,
		37132	=>	19454,
		37133	=>	19451,
		37134	=>	19449,
		37135	=>	19446,
		37136	=>	19443,
		37137	=>	19440,
		37138	=>	19437,
		37139	=>	19434,
		37140	=>	19431,
		37141	=>	19428,
		37142	=>	19426,
		37143	=>	19423,
		37144	=>	19420,
		37145	=>	19417,
		37146	=>	19414,
		37147	=>	19411,
		37148	=>	19408,
		37149	=>	19406,
		37150	=>	19403,
		37151	=>	19400,
		37152	=>	19397,
		37153	=>	19394,
		37154	=>	19391,
		37155	=>	19388,
		37156	=>	19385,
		37157	=>	19383,
		37158	=>	19380,
		37159	=>	19377,
		37160	=>	19374,
		37161	=>	19371,
		37162	=>	19368,
		37163	=>	19365,
		37164	=>	19363,
		37165	=>	19360,
		37166	=>	19357,
		37167	=>	19354,
		37168	=>	19351,
		37169	=>	19348,
		37170	=>	19345,
		37171	=>	19342,
		37172	=>	19340,
		37173	=>	19337,
		37174	=>	19334,
		37175	=>	19331,
		37176	=>	19328,
		37177	=>	19325,
		37178	=>	19322,
		37179	=>	19320,
		37180	=>	19317,
		37181	=>	19314,
		37182	=>	19311,
		37183	=>	19308,
		37184	=>	19305,
		37185	=>	19302,
		37186	=>	19299,
		37187	=>	19297,
		37188	=>	19294,
		37189	=>	19291,
		37190	=>	19288,
		37191	=>	19285,
		37192	=>	19282,
		37193	=>	19279,
		37194	=>	19277,
		37195	=>	19274,
		37196	=>	19271,
		37197	=>	19268,
		37198	=>	19265,
		37199	=>	19262,
		37200	=>	19259,
		37201	=>	19257,
		37202	=>	19254,
		37203	=>	19251,
		37204	=>	19248,
		37205	=>	19245,
		37206	=>	19242,
		37207	=>	19239,
		37208	=>	19236,
		37209	=>	19234,
		37210	=>	19231,
		37211	=>	19228,
		37212	=>	19225,
		37213	=>	19222,
		37214	=>	19219,
		37215	=>	19216,
		37216	=>	19214,
		37217	=>	19211,
		37218	=>	19208,
		37219	=>	19205,
		37220	=>	19202,
		37221	=>	19199,
		37222	=>	19196,
		37223	=>	19194,
		37224	=>	19191,
		37225	=>	19188,
		37226	=>	19185,
		37227	=>	19182,
		37228	=>	19179,
		37229	=>	19176,
		37230	=>	19174,
		37231	=>	19171,
		37232	=>	19168,
		37233	=>	19165,
		37234	=>	19162,
		37235	=>	19159,
		37236	=>	19156,
		37237	=>	19154,
		37238	=>	19151,
		37239	=>	19148,
		37240	=>	19145,
		37241	=>	19142,
		37242	=>	19139,
		37243	=>	19136,
		37244	=>	19134,
		37245	=>	19131,
		37246	=>	19128,
		37247	=>	19125,
		37248	=>	19122,
		37249	=>	19119,
		37250	=>	19116,
		37251	=>	19114,
		37252	=>	19111,
		37253	=>	19108,
		37254	=>	19105,
		37255	=>	19102,
		37256	=>	19099,
		37257	=>	19096,
		37258	=>	19094,
		37259	=>	19091,
		37260	=>	19088,
		37261	=>	19085,
		37262	=>	19082,
		37263	=>	19079,
		37264	=>	19076,
		37265	=>	19074,
		37266	=>	19071,
		37267	=>	19068,
		37268	=>	19065,
		37269	=>	19062,
		37270	=>	19059,
		37271	=>	19056,
		37272	=>	19054,
		37273	=>	19051,
		37274	=>	19048,
		37275	=>	19045,
		37276	=>	19042,
		37277	=>	19039,
		37278	=>	19037,
		37279	=>	19034,
		37280	=>	19031,
		37281	=>	19028,
		37282	=>	19025,
		37283	=>	19022,
		37284	=>	19019,
		37285	=>	19017,
		37286	=>	19014,
		37287	=>	19011,
		37288	=>	19008,
		37289	=>	19005,
		37290	=>	19002,
		37291	=>	18999,
		37292	=>	18997,
		37293	=>	18994,
		37294	=>	18991,
		37295	=>	18988,
		37296	=>	18985,
		37297	=>	18982,
		37298	=>	18979,
		37299	=>	18977,
		37300	=>	18974,
		37301	=>	18971,
		37302	=>	18968,
		37303	=>	18965,
		37304	=>	18962,
		37305	=>	18960,
		37306	=>	18957,
		37307	=>	18954,
		37308	=>	18951,
		37309	=>	18948,
		37310	=>	18945,
		37311	=>	18942,
		37312	=>	18940,
		37313	=>	18937,
		37314	=>	18934,
		37315	=>	18931,
		37316	=>	18928,
		37317	=>	18925,
		37318	=>	18923,
		37319	=>	18920,
		37320	=>	18917,
		37321	=>	18914,
		37322	=>	18911,
		37323	=>	18908,
		37324	=>	18905,
		37325	=>	18903,
		37326	=>	18900,
		37327	=>	18897,
		37328	=>	18894,
		37329	=>	18891,
		37330	=>	18888,
		37331	=>	18886,
		37332	=>	18883,
		37333	=>	18880,
		37334	=>	18877,
		37335	=>	18874,
		37336	=>	18871,
		37337	=>	18868,
		37338	=>	18866,
		37339	=>	18863,
		37340	=>	18860,
		37341	=>	18857,
		37342	=>	18854,
		37343	=>	18851,
		37344	=>	18849,
		37345	=>	18846,
		37346	=>	18843,
		37347	=>	18840,
		37348	=>	18837,
		37349	=>	18834,
		37350	=>	18831,
		37351	=>	18829,
		37352	=>	18826,
		37353	=>	18823,
		37354	=>	18820,
		37355	=>	18817,
		37356	=>	18814,
		37357	=>	18812,
		37358	=>	18809,
		37359	=>	18806,
		37360	=>	18803,
		37361	=>	18800,
		37362	=>	18797,
		37363	=>	18795,
		37364	=>	18792,
		37365	=>	18789,
		37366	=>	18786,
		37367	=>	18783,
		37368	=>	18780,
		37369	=>	18777,
		37370	=>	18775,
		37371	=>	18772,
		37372	=>	18769,
		37373	=>	18766,
		37374	=>	18763,
		37375	=>	18760,
		37376	=>	18758,
		37377	=>	18755,
		37378	=>	18752,
		37379	=>	18749,
		37380	=>	18746,
		37381	=>	18743,
		37382	=>	18741,
		37383	=>	18738,
		37384	=>	18735,
		37385	=>	18732,
		37386	=>	18729,
		37387	=>	18726,
		37388	=>	18724,
		37389	=>	18721,
		37390	=>	18718,
		37391	=>	18715,
		37392	=>	18712,
		37393	=>	18709,
		37394	=>	18706,
		37395	=>	18704,
		37396	=>	18701,
		37397	=>	18698,
		37398	=>	18695,
		37399	=>	18692,
		37400	=>	18689,
		37401	=>	18687,
		37402	=>	18684,
		37403	=>	18681,
		37404	=>	18678,
		37405	=>	18675,
		37406	=>	18672,
		37407	=>	18670,
		37408	=>	18667,
		37409	=>	18664,
		37410	=>	18661,
		37411	=>	18658,
		37412	=>	18655,
		37413	=>	18653,
		37414	=>	18650,
		37415	=>	18647,
		37416	=>	18644,
		37417	=>	18641,
		37418	=>	18638,
		37419	=>	18636,
		37420	=>	18633,
		37421	=>	18630,
		37422	=>	18627,
		37423	=>	18624,
		37424	=>	18621,
		37425	=>	18619,
		37426	=>	18616,
		37427	=>	18613,
		37428	=>	18610,
		37429	=>	18607,
		37430	=>	18604,
		37431	=>	18602,
		37432	=>	18599,
		37433	=>	18596,
		37434	=>	18593,
		37435	=>	18590,
		37436	=>	18587,
		37437	=>	18585,
		37438	=>	18582,
		37439	=>	18579,
		37440	=>	18576,
		37441	=>	18573,
		37442	=>	18570,
		37443	=>	18568,
		37444	=>	18565,
		37445	=>	18562,
		37446	=>	18559,
		37447	=>	18556,
		37448	=>	18553,
		37449	=>	18551,
		37450	=>	18548,
		37451	=>	18545,
		37452	=>	18542,
		37453	=>	18539,
		37454	=>	18536,
		37455	=>	18534,
		37456	=>	18531,
		37457	=>	18528,
		37458	=>	18525,
		37459	=>	18522,
		37460	=>	18519,
		37461	=>	18517,
		37462	=>	18514,
		37463	=>	18511,
		37464	=>	18508,
		37465	=>	18505,
		37466	=>	18503,
		37467	=>	18500,
		37468	=>	18497,
		37469	=>	18494,
		37470	=>	18491,
		37471	=>	18488,
		37472	=>	18486,
		37473	=>	18483,
		37474	=>	18480,
		37475	=>	18477,
		37476	=>	18474,
		37477	=>	18471,
		37478	=>	18469,
		37479	=>	18466,
		37480	=>	18463,
		37481	=>	18460,
		37482	=>	18457,
		37483	=>	18454,
		37484	=>	18452,
		37485	=>	18449,
		37486	=>	18446,
		37487	=>	18443,
		37488	=>	18440,
		37489	=>	18438,
		37490	=>	18435,
		37491	=>	18432,
		37492	=>	18429,
		37493	=>	18426,
		37494	=>	18423,
		37495	=>	18421,
		37496	=>	18418,
		37497	=>	18415,
		37498	=>	18412,
		37499	=>	18409,
		37500	=>	18406,
		37501	=>	18404,
		37502	=>	18401,
		37503	=>	18398,
		37504	=>	18395,
		37505	=>	18392,
		37506	=>	18389,
		37507	=>	18387,
		37508	=>	18384,
		37509	=>	18381,
		37510	=>	18378,
		37511	=>	18375,
		37512	=>	18373,
		37513	=>	18370,
		37514	=>	18367,
		37515	=>	18364,
		37516	=>	18361,
		37517	=>	18358,
		37518	=>	18356,
		37519	=>	18353,
		37520	=>	18350,
		37521	=>	18347,
		37522	=>	18344,
		37523	=>	18342,
		37524	=>	18339,
		37525	=>	18336,
		37526	=>	18333,
		37527	=>	18330,
		37528	=>	18327,
		37529	=>	18325,
		37530	=>	18322,
		37531	=>	18319,
		37532	=>	18316,
		37533	=>	18313,
		37534	=>	18311,
		37535	=>	18308,
		37536	=>	18305,
		37537	=>	18302,
		37538	=>	18299,
		37539	=>	18296,
		37540	=>	18294,
		37541	=>	18291,
		37542	=>	18288,
		37543	=>	18285,
		37544	=>	18282,
		37545	=>	18280,
		37546	=>	18277,
		37547	=>	18274,
		37548	=>	18271,
		37549	=>	18268,
		37550	=>	18265,
		37551	=>	18263,
		37552	=>	18260,
		37553	=>	18257,
		37554	=>	18254,
		37555	=>	18251,
		37556	=>	18249,
		37557	=>	18246,
		37558	=>	18243,
		37559	=>	18240,
		37560	=>	18237,
		37561	=>	18234,
		37562	=>	18232,
		37563	=>	18229,
		37564	=>	18226,
		37565	=>	18223,
		37566	=>	18220,
		37567	=>	18218,
		37568	=>	18215,
		37569	=>	18212,
		37570	=>	18209,
		37571	=>	18206,
		37572	=>	18203,
		37573	=>	18201,
		37574	=>	18198,
		37575	=>	18195,
		37576	=>	18192,
		37577	=>	18189,
		37578	=>	18187,
		37579	=>	18184,
		37580	=>	18181,
		37581	=>	18178,
		37582	=>	18175,
		37583	=>	18173,
		37584	=>	18170,
		37585	=>	18167,
		37586	=>	18164,
		37587	=>	18161,
		37588	=>	18158,
		37589	=>	18156,
		37590	=>	18153,
		37591	=>	18150,
		37592	=>	18147,
		37593	=>	18144,
		37594	=>	18142,
		37595	=>	18139,
		37596	=>	18136,
		37597	=>	18133,
		37598	=>	18130,
		37599	=>	18128,
		37600	=>	18125,
		37601	=>	18122,
		37602	=>	18119,
		37603	=>	18116,
		37604	=>	18113,
		37605	=>	18111,
		37606	=>	18108,
		37607	=>	18105,
		37608	=>	18102,
		37609	=>	18099,
		37610	=>	18097,
		37611	=>	18094,
		37612	=>	18091,
		37613	=>	18088,
		37614	=>	18085,
		37615	=>	18083,
		37616	=>	18080,
		37617	=>	18077,
		37618	=>	18074,
		37619	=>	18071,
		37620	=>	18069,
		37621	=>	18066,
		37622	=>	18063,
		37623	=>	18060,
		37624	=>	18057,
		37625	=>	18055,
		37626	=>	18052,
		37627	=>	18049,
		37628	=>	18046,
		37629	=>	18043,
		37630	=>	18040,
		37631	=>	18038,
		37632	=>	18035,
		37633	=>	18032,
		37634	=>	18029,
		37635	=>	18026,
		37636	=>	18024,
		37637	=>	18021,
		37638	=>	18018,
		37639	=>	18015,
		37640	=>	18012,
		37641	=>	18010,
		37642	=>	18007,
		37643	=>	18004,
		37644	=>	18001,
		37645	=>	17998,
		37646	=>	17996,
		37647	=>	17993,
		37648	=>	17990,
		37649	=>	17987,
		37650	=>	17984,
		37651	=>	17982,
		37652	=>	17979,
		37653	=>	17976,
		37654	=>	17973,
		37655	=>	17970,
		37656	=>	17968,
		37657	=>	17965,
		37658	=>	17962,
		37659	=>	17959,
		37660	=>	17956,
		37661	=>	17954,
		37662	=>	17951,
		37663	=>	17948,
		37664	=>	17945,
		37665	=>	17942,
		37666	=>	17940,
		37667	=>	17937,
		37668	=>	17934,
		37669	=>	17931,
		37670	=>	17928,
		37671	=>	17926,
		37672	=>	17923,
		37673	=>	17920,
		37674	=>	17917,
		37675	=>	17914,
		37676	=>	17912,
		37677	=>	17909,
		37678	=>	17906,
		37679	=>	17903,
		37680	=>	17900,
		37681	=>	17898,
		37682	=>	17895,
		37683	=>	17892,
		37684	=>	17889,
		37685	=>	17886,
		37686	=>	17884,
		37687	=>	17881,
		37688	=>	17878,
		37689	=>	17875,
		37690	=>	17872,
		37691	=>	17870,
		37692	=>	17867,
		37693	=>	17864,
		37694	=>	17861,
		37695	=>	17858,
		37696	=>	17856,
		37697	=>	17853,
		37698	=>	17850,
		37699	=>	17847,
		37700	=>	17844,
		37701	=>	17842,
		37702	=>	17839,
		37703	=>	17836,
		37704	=>	17833,
		37705	=>	17830,
		37706	=>	17828,
		37707	=>	17825,
		37708	=>	17822,
		37709	=>	17819,
		37710	=>	17816,
		37711	=>	17814,
		37712	=>	17811,
		37713	=>	17808,
		37714	=>	17805,
		37715	=>	17802,
		37716	=>	17800,
		37717	=>	17797,
		37718	=>	17794,
		37719	=>	17791,
		37720	=>	17788,
		37721	=>	17786,
		37722	=>	17783,
		37723	=>	17780,
		37724	=>	17777,
		37725	=>	17774,
		37726	=>	17772,
		37727	=>	17769,
		37728	=>	17766,
		37729	=>	17763,
		37730	=>	17761,
		37731	=>	17758,
		37732	=>	17755,
		37733	=>	17752,
		37734	=>	17749,
		37735	=>	17747,
		37736	=>	17744,
		37737	=>	17741,
		37738	=>	17738,
		37739	=>	17735,
		37740	=>	17733,
		37741	=>	17730,
		37742	=>	17727,
		37743	=>	17724,
		37744	=>	17721,
		37745	=>	17719,
		37746	=>	17716,
		37747	=>	17713,
		37748	=>	17710,
		37749	=>	17707,
		37750	=>	17705,
		37751	=>	17702,
		37752	=>	17699,
		37753	=>	17696,
		37754	=>	17694,
		37755	=>	17691,
		37756	=>	17688,
		37757	=>	17685,
		37758	=>	17682,
		37759	=>	17680,
		37760	=>	17677,
		37761	=>	17674,
		37762	=>	17671,
		37763	=>	17668,
		37764	=>	17666,
		37765	=>	17663,
		37766	=>	17660,
		37767	=>	17657,
		37768	=>	17654,
		37769	=>	17652,
		37770	=>	17649,
		37771	=>	17646,
		37772	=>	17643,
		37773	=>	17641,
		37774	=>	17638,
		37775	=>	17635,
		37776	=>	17632,
		37777	=>	17629,
		37778	=>	17627,
		37779	=>	17624,
		37780	=>	17621,
		37781	=>	17618,
		37782	=>	17615,
		37783	=>	17613,
		37784	=>	17610,
		37785	=>	17607,
		37786	=>	17604,
		37787	=>	17602,
		37788	=>	17599,
		37789	=>	17596,
		37790	=>	17593,
		37791	=>	17590,
		37792	=>	17588,
		37793	=>	17585,
		37794	=>	17582,
		37795	=>	17579,
		37796	=>	17576,
		37797	=>	17574,
		37798	=>	17571,
		37799	=>	17568,
		37800	=>	17565,
		37801	=>	17563,
		37802	=>	17560,
		37803	=>	17557,
		37804	=>	17554,
		37805	=>	17551,
		37806	=>	17549,
		37807	=>	17546,
		37808	=>	17543,
		37809	=>	17540,
		37810	=>	17538,
		37811	=>	17535,
		37812	=>	17532,
		37813	=>	17529,
		37814	=>	17526,
		37815	=>	17524,
		37816	=>	17521,
		37817	=>	17518,
		37818	=>	17515,
		37819	=>	17513,
		37820	=>	17510,
		37821	=>	17507,
		37822	=>	17504,
		37823	=>	17501,
		37824	=>	17499,
		37825	=>	17496,
		37826	=>	17493,
		37827	=>	17490,
		37828	=>	17487,
		37829	=>	17485,
		37830	=>	17482,
		37831	=>	17479,
		37832	=>	17476,
		37833	=>	17474,
		37834	=>	17471,
		37835	=>	17468,
		37836	=>	17465,
		37837	=>	17462,
		37838	=>	17460,
		37839	=>	17457,
		37840	=>	17454,
		37841	=>	17451,
		37842	=>	17449,
		37843	=>	17446,
		37844	=>	17443,
		37845	=>	17440,
		37846	=>	17437,
		37847	=>	17435,
		37848	=>	17432,
		37849	=>	17429,
		37850	=>	17426,
		37851	=>	17424,
		37852	=>	17421,
		37853	=>	17418,
		37854	=>	17415,
		37855	=>	17413,
		37856	=>	17410,
		37857	=>	17407,
		37858	=>	17404,
		37859	=>	17401,
		37860	=>	17399,
		37861	=>	17396,
		37862	=>	17393,
		37863	=>	17390,
		37864	=>	17388,
		37865	=>	17385,
		37866	=>	17382,
		37867	=>	17379,
		37868	=>	17376,
		37869	=>	17374,
		37870	=>	17371,
		37871	=>	17368,
		37872	=>	17365,
		37873	=>	17363,
		37874	=>	17360,
		37875	=>	17357,
		37876	=>	17354,
		37877	=>	17351,
		37878	=>	17349,
		37879	=>	17346,
		37880	=>	17343,
		37881	=>	17340,
		37882	=>	17338,
		37883	=>	17335,
		37884	=>	17332,
		37885	=>	17329,
		37886	=>	17327,
		37887	=>	17324,
		37888	=>	17321,
		37889	=>	17318,
		37890	=>	17315,
		37891	=>	17313,
		37892	=>	17310,
		37893	=>	17307,
		37894	=>	17304,
		37895	=>	17302,
		37896	=>	17299,
		37897	=>	17296,
		37898	=>	17293,
		37899	=>	17291,
		37900	=>	17288,
		37901	=>	17285,
		37902	=>	17282,
		37903	=>	17279,
		37904	=>	17277,
		37905	=>	17274,
		37906	=>	17271,
		37907	=>	17268,
		37908	=>	17266,
		37909	=>	17263,
		37910	=>	17260,
		37911	=>	17257,
		37912	=>	17255,
		37913	=>	17252,
		37914	=>	17249,
		37915	=>	17246,
		37916	=>	17243,
		37917	=>	17241,
		37918	=>	17238,
		37919	=>	17235,
		37920	=>	17232,
		37921	=>	17230,
		37922	=>	17227,
		37923	=>	17224,
		37924	=>	17221,
		37925	=>	17219,
		37926	=>	17216,
		37927	=>	17213,
		37928	=>	17210,
		37929	=>	17208,
		37930	=>	17205,
		37931	=>	17202,
		37932	=>	17199,
		37933	=>	17196,
		37934	=>	17194,
		37935	=>	17191,
		37936	=>	17188,
		37937	=>	17185,
		37938	=>	17183,
		37939	=>	17180,
		37940	=>	17177,
		37941	=>	17174,
		37942	=>	17172,
		37943	=>	17169,
		37944	=>	17166,
		37945	=>	17163,
		37946	=>	17161,
		37947	=>	17158,
		37948	=>	17155,
		37949	=>	17152,
		37950	=>	17150,
		37951	=>	17147,
		37952	=>	17144,
		37953	=>	17141,
		37954	=>	17138,
		37955	=>	17136,
		37956	=>	17133,
		37957	=>	17130,
		37958	=>	17127,
		37959	=>	17125,
		37960	=>	17122,
		37961	=>	17119,
		37962	=>	17116,
		37963	=>	17114,
		37964	=>	17111,
		37965	=>	17108,
		37966	=>	17105,
		37967	=>	17103,
		37968	=>	17100,
		37969	=>	17097,
		37970	=>	17094,
		37971	=>	17092,
		37972	=>	17089,
		37973	=>	17086,
		37974	=>	17083,
		37975	=>	17081,
		37976	=>	17078,
		37977	=>	17075,
		37978	=>	17072,
		37979	=>	17069,
		37980	=>	17067,
		37981	=>	17064,
		37982	=>	17061,
		37983	=>	17058,
		37984	=>	17056,
		37985	=>	17053,
		37986	=>	17050,
		37987	=>	17047,
		37988	=>	17045,
		37989	=>	17042,
		37990	=>	17039,
		37991	=>	17036,
		37992	=>	17034,
		37993	=>	17031,
		37994	=>	17028,
		37995	=>	17025,
		37996	=>	17023,
		37997	=>	17020,
		37998	=>	17017,
		37999	=>	17014,
		38000	=>	17012,
		38001	=>	17009,
		38002	=>	17006,
		38003	=>	17003,
		38004	=>	17001,
		38005	=>	16998,
		38006	=>	16995,
		38007	=>	16992,
		38008	=>	16990,
		38009	=>	16987,
		38010	=>	16984,
		38011	=>	16981,
		38012	=>	16979,
		38013	=>	16976,
		38014	=>	16973,
		38015	=>	16970,
		38016	=>	16968,
		38017	=>	16965,
		38018	=>	16962,
		38019	=>	16959,
		38020	=>	16957,
		38021	=>	16954,
		38022	=>	16951,
		38023	=>	16948,
		38024	=>	16946,
		38025	=>	16943,
		38026	=>	16940,
		38027	=>	16937,
		38028	=>	16935,
		38029	=>	16932,
		38030	=>	16929,
		38031	=>	16926,
		38032	=>	16924,
		38033	=>	16921,
		38034	=>	16918,
		38035	=>	16915,
		38036	=>	16913,
		38037	=>	16910,
		38038	=>	16907,
		38039	=>	16904,
		38040	=>	16902,
		38041	=>	16899,
		38042	=>	16896,
		38043	=>	16893,
		38044	=>	16891,
		38045	=>	16888,
		38046	=>	16885,
		38047	=>	16882,
		38048	=>	16880,
		38049	=>	16877,
		38050	=>	16874,
		38051	=>	16871,
		38052	=>	16869,
		38053	=>	16866,
		38054	=>	16863,
		38055	=>	16860,
		38056	=>	16858,
		38057	=>	16855,
		38058	=>	16852,
		38059	=>	16849,
		38060	=>	16847,
		38061	=>	16844,
		38062	=>	16841,
		38063	=>	16838,
		38064	=>	16836,
		38065	=>	16833,
		38066	=>	16830,
		38067	=>	16827,
		38068	=>	16825,
		38069	=>	16822,
		38070	=>	16819,
		38071	=>	16816,
		38072	=>	16814,
		38073	=>	16811,
		38074	=>	16808,
		38075	=>	16805,
		38076	=>	16803,
		38077	=>	16800,
		38078	=>	16797,
		38079	=>	16794,
		38080	=>	16792,
		38081	=>	16789,
		38082	=>	16786,
		38083	=>	16783,
		38084	=>	16781,
		38085	=>	16778,
		38086	=>	16775,
		38087	=>	16773,
		38088	=>	16770,
		38089	=>	16767,
		38090	=>	16764,
		38091	=>	16762,
		38092	=>	16759,
		38093	=>	16756,
		38094	=>	16753,
		38095	=>	16751,
		38096	=>	16748,
		38097	=>	16745,
		38098	=>	16742,
		38099	=>	16740,
		38100	=>	16737,
		38101	=>	16734,
		38102	=>	16731,
		38103	=>	16729,
		38104	=>	16726,
		38105	=>	16723,
		38106	=>	16720,
		38107	=>	16718,
		38108	=>	16715,
		38109	=>	16712,
		38110	=>	16709,
		38111	=>	16707,
		38112	=>	16704,
		38113	=>	16701,
		38114	=>	16699,
		38115	=>	16696,
		38116	=>	16693,
		38117	=>	16690,
		38118	=>	16688,
		38119	=>	16685,
		38120	=>	16682,
		38121	=>	16679,
		38122	=>	16677,
		38123	=>	16674,
		38124	=>	16671,
		38125	=>	16668,
		38126	=>	16666,
		38127	=>	16663,
		38128	=>	16660,
		38129	=>	16657,
		38130	=>	16655,
		38131	=>	16652,
		38132	=>	16649,
		38133	=>	16647,
		38134	=>	16644,
		38135	=>	16641,
		38136	=>	16638,
		38137	=>	16636,
		38138	=>	16633,
		38139	=>	16630,
		38140	=>	16627,
		38141	=>	16625,
		38142	=>	16622,
		38143	=>	16619,
		38144	=>	16616,
		38145	=>	16614,
		38146	=>	16611,
		38147	=>	16608,
		38148	=>	16606,
		38149	=>	16603,
		38150	=>	16600,
		38151	=>	16597,
		38152	=>	16595,
		38153	=>	16592,
		38154	=>	16589,
		38155	=>	16586,
		38156	=>	16584,
		38157	=>	16581,
		38158	=>	16578,
		38159	=>	16575,
		38160	=>	16573,
		38161	=>	16570,
		38162	=>	16567,
		38163	=>	16565,
		38164	=>	16562,
		38165	=>	16559,
		38166	=>	16556,
		38167	=>	16554,
		38168	=>	16551,
		38169	=>	16548,
		38170	=>	16545,
		38171	=>	16543,
		38172	=>	16540,
		38173	=>	16537,
		38174	=>	16535,
		38175	=>	16532,
		38176	=>	16529,
		38177	=>	16526,
		38178	=>	16524,
		38179	=>	16521,
		38180	=>	16518,
		38181	=>	16515,
		38182	=>	16513,
		38183	=>	16510,
		38184	=>	16507,
		38185	=>	16505,
		38186	=>	16502,
		38187	=>	16499,
		38188	=>	16496,
		38189	=>	16494,
		38190	=>	16491,
		38191	=>	16488,
		38192	=>	16485,
		38193	=>	16483,
		38194	=>	16480,
		38195	=>	16477,
		38196	=>	16475,
		38197	=>	16472,
		38198	=>	16469,
		38199	=>	16466,
		38200	=>	16464,
		38201	=>	16461,
		38202	=>	16458,
		38203	=>	16455,
		38204	=>	16453,
		38205	=>	16450,
		38206	=>	16447,
		38207	=>	16445,
		38208	=>	16442,
		38209	=>	16439,
		38210	=>	16436,
		38211	=>	16434,
		38212	=>	16431,
		38213	=>	16428,
		38214	=>	16425,
		38215	=>	16423,
		38216	=>	16420,
		38217	=>	16417,
		38218	=>	16415,
		38219	=>	16412,
		38220	=>	16409,
		38221	=>	16406,
		38222	=>	16404,
		38223	=>	16401,
		38224	=>	16398,
		38225	=>	16396,
		38226	=>	16393,
		38227	=>	16390,
		38228	=>	16387,
		38229	=>	16385,
		38230	=>	16382,
		38231	=>	16379,
		38232	=>	16376,
		38233	=>	16374,
		38234	=>	16371,
		38235	=>	16368,
		38236	=>	16366,
		38237	=>	16363,
		38238	=>	16360,
		38239	=>	16357,
		38240	=>	16355,
		38241	=>	16352,
		38242	=>	16349,
		38243	=>	16347,
		38244	=>	16344,
		38245	=>	16341,
		38246	=>	16338,
		38247	=>	16336,
		38248	=>	16333,
		38249	=>	16330,
		38250	=>	16328,
		38251	=>	16325,
		38252	=>	16322,
		38253	=>	16319,
		38254	=>	16317,
		38255	=>	16314,
		38256	=>	16311,
		38257	=>	16309,
		38258	=>	16306,
		38259	=>	16303,
		38260	=>	16300,
		38261	=>	16298,
		38262	=>	16295,
		38263	=>	16292,
		38264	=>	16290,
		38265	=>	16287,
		38266	=>	16284,
		38267	=>	16281,
		38268	=>	16279,
		38269	=>	16276,
		38270	=>	16273,
		38271	=>	16271,
		38272	=>	16268,
		38273	=>	16265,
		38274	=>	16262,
		38275	=>	16260,
		38276	=>	16257,
		38277	=>	16254,
		38278	=>	16252,
		38279	=>	16249,
		38280	=>	16246,
		38281	=>	16243,
		38282	=>	16241,
		38283	=>	16238,
		38284	=>	16235,
		38285	=>	16233,
		38286	=>	16230,
		38287	=>	16227,
		38288	=>	16224,
		38289	=>	16222,
		38290	=>	16219,
		38291	=>	16216,
		38292	=>	16214,
		38293	=>	16211,
		38294	=>	16208,
		38295	=>	16205,
		38296	=>	16203,
		38297	=>	16200,
		38298	=>	16197,
		38299	=>	16195,
		38300	=>	16192,
		38301	=>	16189,
		38302	=>	16186,
		38303	=>	16184,
		38304	=>	16181,
		38305	=>	16178,
		38306	=>	16176,
		38307	=>	16173,
		38308	=>	16170,
		38309	=>	16167,
		38310	=>	16165,
		38311	=>	16162,
		38312	=>	16159,
		38313	=>	16157,
		38314	=>	16154,
		38315	=>	16151,
		38316	=>	16149,
		38317	=>	16146,
		38318	=>	16143,
		38319	=>	16140,
		38320	=>	16138,
		38321	=>	16135,
		38322	=>	16132,
		38323	=>	16130,
		38324	=>	16127,
		38325	=>	16124,
		38326	=>	16121,
		38327	=>	16119,
		38328	=>	16116,
		38329	=>	16113,
		38330	=>	16111,
		38331	=>	16108,
		38332	=>	16105,
		38333	=>	16103,
		38334	=>	16100,
		38335	=>	16097,
		38336	=>	16094,
		38337	=>	16092,
		38338	=>	16089,
		38339	=>	16086,
		38340	=>	16084,
		38341	=>	16081,
		38342	=>	16078,
		38343	=>	16075,
		38344	=>	16073,
		38345	=>	16070,
		38346	=>	16067,
		38347	=>	16065,
		38348	=>	16062,
		38349	=>	16059,
		38350	=>	16057,
		38351	=>	16054,
		38352	=>	16051,
		38353	=>	16048,
		38354	=>	16046,
		38355	=>	16043,
		38356	=>	16040,
		38357	=>	16038,
		38358	=>	16035,
		38359	=>	16032,
		38360	=>	16030,
		38361	=>	16027,
		38362	=>	16024,
		38363	=>	16021,
		38364	=>	16019,
		38365	=>	16016,
		38366	=>	16013,
		38367	=>	16011,
		38368	=>	16008,
		38369	=>	16005,
		38370	=>	16003,
		38371	=>	16000,
		38372	=>	15997,
		38373	=>	15994,
		38374	=>	15992,
		38375	=>	15989,
		38376	=>	15986,
		38377	=>	15984,
		38378	=>	15981,
		38379	=>	15978,
		38380	=>	15976,
		38381	=>	15973,
		38382	=>	15970,
		38383	=>	15967,
		38384	=>	15965,
		38385	=>	15962,
		38386	=>	15959,
		38387	=>	15957,
		38388	=>	15954,
		38389	=>	15951,
		38390	=>	15949,
		38391	=>	15946,
		38392	=>	15943,
		38393	=>	15941,
		38394	=>	15938,
		38395	=>	15935,
		38396	=>	15932,
		38397	=>	15930,
		38398	=>	15927,
		38399	=>	15924,
		38400	=>	15922,
		38401	=>	15919,
		38402	=>	15916,
		38403	=>	15914,
		38404	=>	15911,
		38405	=>	15908,
		38406	=>	15905,
		38407	=>	15903,
		38408	=>	15900,
		38409	=>	15897,
		38410	=>	15895,
		38411	=>	15892,
		38412	=>	15889,
		38413	=>	15887,
		38414	=>	15884,
		38415	=>	15881,
		38416	=>	15879,
		38417	=>	15876,
		38418	=>	15873,
		38419	=>	15870,
		38420	=>	15868,
		38421	=>	15865,
		38422	=>	15862,
		38423	=>	15860,
		38424	=>	15857,
		38425	=>	15854,
		38426	=>	15852,
		38427	=>	15849,
		38428	=>	15846,
		38429	=>	15844,
		38430	=>	15841,
		38431	=>	15838,
		38432	=>	15835,
		38433	=>	15833,
		38434	=>	15830,
		38435	=>	15827,
		38436	=>	15825,
		38437	=>	15822,
		38438	=>	15819,
		38439	=>	15817,
		38440	=>	15814,
		38441	=>	15811,
		38442	=>	15809,
		38443	=>	15806,
		38444	=>	15803,
		38445	=>	15801,
		38446	=>	15798,
		38447	=>	15795,
		38448	=>	15792,
		38449	=>	15790,
		38450	=>	15787,
		38451	=>	15784,
		38452	=>	15782,
		38453	=>	15779,
		38454	=>	15776,
		38455	=>	15774,
		38456	=>	15771,
		38457	=>	15768,
		38458	=>	15766,
		38459	=>	15763,
		38460	=>	15760,
		38461	=>	15758,
		38462	=>	15755,
		38463	=>	15752,
		38464	=>	15750,
		38465	=>	15747,
		38466	=>	15744,
		38467	=>	15741,
		38468	=>	15739,
		38469	=>	15736,
		38470	=>	15733,
		38471	=>	15731,
		38472	=>	15728,
		38473	=>	15725,
		38474	=>	15723,
		38475	=>	15720,
		38476	=>	15717,
		38477	=>	15715,
		38478	=>	15712,
		38479	=>	15709,
		38480	=>	15707,
		38481	=>	15704,
		38482	=>	15701,
		38483	=>	15699,
		38484	=>	15696,
		38485	=>	15693,
		38486	=>	15690,
		38487	=>	15688,
		38488	=>	15685,
		38489	=>	15682,
		38490	=>	15680,
		38491	=>	15677,
		38492	=>	15674,
		38493	=>	15672,
		38494	=>	15669,
		38495	=>	15666,
		38496	=>	15664,
		38497	=>	15661,
		38498	=>	15658,
		38499	=>	15656,
		38500	=>	15653,
		38501	=>	15650,
		38502	=>	15648,
		38503	=>	15645,
		38504	=>	15642,
		38505	=>	15640,
		38506	=>	15637,
		38507	=>	15634,
		38508	=>	15632,
		38509	=>	15629,
		38510	=>	15626,
		38511	=>	15623,
		38512	=>	15621,
		38513	=>	15618,
		38514	=>	15615,
		38515	=>	15613,
		38516	=>	15610,
		38517	=>	15607,
		38518	=>	15605,
		38519	=>	15602,
		38520	=>	15599,
		38521	=>	15597,
		38522	=>	15594,
		38523	=>	15591,
		38524	=>	15589,
		38525	=>	15586,
		38526	=>	15583,
		38527	=>	15581,
		38528	=>	15578,
		38529	=>	15575,
		38530	=>	15573,
		38531	=>	15570,
		38532	=>	15567,
		38533	=>	15565,
		38534	=>	15562,
		38535	=>	15559,
		38536	=>	15557,
		38537	=>	15554,
		38538	=>	15551,
		38539	=>	15549,
		38540	=>	15546,
		38541	=>	15543,
		38542	=>	15541,
		38543	=>	15538,
		38544	=>	15535,
		38545	=>	15533,
		38546	=>	15530,
		38547	=>	15527,
		38548	=>	15525,
		38549	=>	15522,
		38550	=>	15519,
		38551	=>	15517,
		38552	=>	15514,
		38553	=>	15511,
		38554	=>	15509,
		38555	=>	15506,
		38556	=>	15503,
		38557	=>	15501,
		38558	=>	15498,
		38559	=>	15495,
		38560	=>	15493,
		38561	=>	15490,
		38562	=>	15487,
		38563	=>	15484,
		38564	=>	15482,
		38565	=>	15479,
		38566	=>	15476,
		38567	=>	15474,
		38568	=>	15471,
		38569	=>	15468,
		38570	=>	15466,
		38571	=>	15463,
		38572	=>	15460,
		38573	=>	15458,
		38574	=>	15455,
		38575	=>	15452,
		38576	=>	15450,
		38577	=>	15447,
		38578	=>	15444,
		38579	=>	15442,
		38580	=>	15439,
		38581	=>	15436,
		38582	=>	15434,
		38583	=>	15431,
		38584	=>	15428,
		38585	=>	15426,
		38586	=>	15423,
		38587	=>	15420,
		38588	=>	15418,
		38589	=>	15415,
		38590	=>	15412,
		38591	=>	15410,
		38592	=>	15407,
		38593	=>	15404,
		38594	=>	15402,
		38595	=>	15399,
		38596	=>	15397,
		38597	=>	15394,
		38598	=>	15391,
		38599	=>	15389,
		38600	=>	15386,
		38601	=>	15383,
		38602	=>	15381,
		38603	=>	15378,
		38604	=>	15375,
		38605	=>	15373,
		38606	=>	15370,
		38607	=>	15367,
		38608	=>	15365,
		38609	=>	15362,
		38610	=>	15359,
		38611	=>	15357,
		38612	=>	15354,
		38613	=>	15351,
		38614	=>	15349,
		38615	=>	15346,
		38616	=>	15343,
		38617	=>	15341,
		38618	=>	15338,
		38619	=>	15335,
		38620	=>	15333,
		38621	=>	15330,
		38622	=>	15327,
		38623	=>	15325,
		38624	=>	15322,
		38625	=>	15319,
		38626	=>	15317,
		38627	=>	15314,
		38628	=>	15311,
		38629	=>	15309,
		38630	=>	15306,
		38631	=>	15303,
		38632	=>	15301,
		38633	=>	15298,
		38634	=>	15295,
		38635	=>	15293,
		38636	=>	15290,
		38637	=>	15287,
		38638	=>	15285,
		38639	=>	15282,
		38640	=>	15279,
		38641	=>	15277,
		38642	=>	15274,
		38643	=>	15271,
		38644	=>	15269,
		38645	=>	15266,
		38646	=>	15264,
		38647	=>	15261,
		38648	=>	15258,
		38649	=>	15256,
		38650	=>	15253,
		38651	=>	15250,
		38652	=>	15248,
		38653	=>	15245,
		38654	=>	15242,
		38655	=>	15240,
		38656	=>	15237,
		38657	=>	15234,
		38658	=>	15232,
		38659	=>	15229,
		38660	=>	15226,
		38661	=>	15224,
		38662	=>	15221,
		38663	=>	15218,
		38664	=>	15216,
		38665	=>	15213,
		38666	=>	15210,
		38667	=>	15208,
		38668	=>	15205,
		38669	=>	15202,
		38670	=>	15200,
		38671	=>	15197,
		38672	=>	15195,
		38673	=>	15192,
		38674	=>	15189,
		38675	=>	15187,
		38676	=>	15184,
		38677	=>	15181,
		38678	=>	15179,
		38679	=>	15176,
		38680	=>	15173,
		38681	=>	15171,
		38682	=>	15168,
		38683	=>	15165,
		38684	=>	15163,
		38685	=>	15160,
		38686	=>	15157,
		38687	=>	15155,
		38688	=>	15152,
		38689	=>	15149,
		38690	=>	15147,
		38691	=>	15144,
		38692	=>	15142,
		38693	=>	15139,
		38694	=>	15136,
		38695	=>	15134,
		38696	=>	15131,
		38697	=>	15128,
		38698	=>	15126,
		38699	=>	15123,
		38700	=>	15120,
		38701	=>	15118,
		38702	=>	15115,
		38703	=>	15112,
		38704	=>	15110,
		38705	=>	15107,
		38706	=>	15104,
		38707	=>	15102,
		38708	=>	15099,
		38709	=>	15097,
		38710	=>	15094,
		38711	=>	15091,
		38712	=>	15089,
		38713	=>	15086,
		38714	=>	15083,
		38715	=>	15081,
		38716	=>	15078,
		38717	=>	15075,
		38718	=>	15073,
		38719	=>	15070,
		38720	=>	15067,
		38721	=>	15065,
		38722	=>	15062,
		38723	=>	15060,
		38724	=>	15057,
		38725	=>	15054,
		38726	=>	15052,
		38727	=>	15049,
		38728	=>	15046,
		38729	=>	15044,
		38730	=>	15041,
		38731	=>	15038,
		38732	=>	15036,
		38733	=>	15033,
		38734	=>	15030,
		38735	=>	15028,
		38736	=>	15025,
		38737	=>	15023,
		38738	=>	15020,
		38739	=>	15017,
		38740	=>	15015,
		38741	=>	15012,
		38742	=>	15009,
		38743	=>	15007,
		38744	=>	15004,
		38745	=>	15001,
		38746	=>	14999,
		38747	=>	14996,
		38748	=>	14993,
		38749	=>	14991,
		38750	=>	14988,
		38751	=>	14986,
		38752	=>	14983,
		38753	=>	14980,
		38754	=>	14978,
		38755	=>	14975,
		38756	=>	14972,
		38757	=>	14970,
		38758	=>	14967,
		38759	=>	14964,
		38760	=>	14962,
		38761	=>	14959,
		38762	=>	14957,
		38763	=>	14954,
		38764	=>	14951,
		38765	=>	14949,
		38766	=>	14946,
		38767	=>	14943,
		38768	=>	14941,
		38769	=>	14938,
		38770	=>	14935,
		38771	=>	14933,
		38772	=>	14930,
		38773	=>	14928,
		38774	=>	14925,
		38775	=>	14922,
		38776	=>	14920,
		38777	=>	14917,
		38778	=>	14914,
		38779	=>	14912,
		38780	=>	14909,
		38781	=>	14906,
		38782	=>	14904,
		38783	=>	14901,
		38784	=>	14899,
		38785	=>	14896,
		38786	=>	14893,
		38787	=>	14891,
		38788	=>	14888,
		38789	=>	14885,
		38790	=>	14883,
		38791	=>	14880,
		38792	=>	14878,
		38793	=>	14875,
		38794	=>	14872,
		38795	=>	14870,
		38796	=>	14867,
		38797	=>	14864,
		38798	=>	14862,
		38799	=>	14859,
		38800	=>	14856,
		38801	=>	14854,
		38802	=>	14851,
		38803	=>	14849,
		38804	=>	14846,
		38805	=>	14843,
		38806	=>	14841,
		38807	=>	14838,
		38808	=>	14835,
		38809	=>	14833,
		38810	=>	14830,
		38811	=>	14828,
		38812	=>	14825,
		38813	=>	14822,
		38814	=>	14820,
		38815	=>	14817,
		38816	=>	14814,
		38817	=>	14812,
		38818	=>	14809,
		38819	=>	14806,
		38820	=>	14804,
		38821	=>	14801,
		38822	=>	14799,
		38823	=>	14796,
		38824	=>	14793,
		38825	=>	14791,
		38826	=>	14788,
		38827	=>	14785,
		38828	=>	14783,
		38829	=>	14780,
		38830	=>	14778,
		38831	=>	14775,
		38832	=>	14772,
		38833	=>	14770,
		38834	=>	14767,
		38835	=>	14764,
		38836	=>	14762,
		38837	=>	14759,
		38838	=>	14757,
		38839	=>	14754,
		38840	=>	14751,
		38841	=>	14749,
		38842	=>	14746,
		38843	=>	14743,
		38844	=>	14741,
		38845	=>	14738,
		38846	=>	14736,
		38847	=>	14733,
		38848	=>	14730,
		38849	=>	14728,
		38850	=>	14725,
		38851	=>	14723,
		38852	=>	14720,
		38853	=>	14717,
		38854	=>	14715,
		38855	=>	14712,
		38856	=>	14709,
		38857	=>	14707,
		38858	=>	14704,
		38859	=>	14702,
		38860	=>	14699,
		38861	=>	14696,
		38862	=>	14694,
		38863	=>	14691,
		38864	=>	14688,
		38865	=>	14686,
		38866	=>	14683,
		38867	=>	14681,
		38868	=>	14678,
		38869	=>	14675,
		38870	=>	14673,
		38871	=>	14670,
		38872	=>	14667,
		38873	=>	14665,
		38874	=>	14662,
		38875	=>	14660,
		38876	=>	14657,
		38877	=>	14654,
		38878	=>	14652,
		38879	=>	14649,
		38880	=>	14647,
		38881	=>	14644,
		38882	=>	14641,
		38883	=>	14639,
		38884	=>	14636,
		38885	=>	14633,
		38886	=>	14631,
		38887	=>	14628,
		38888	=>	14626,
		38889	=>	14623,
		38890	=>	14620,
		38891	=>	14618,
		38892	=>	14615,
		38893	=>	14613,
		38894	=>	14610,
		38895	=>	14607,
		38896	=>	14605,
		38897	=>	14602,
		38898	=>	14599,
		38899	=>	14597,
		38900	=>	14594,
		38901	=>	14592,
		38902	=>	14589,
		38903	=>	14586,
		38904	=>	14584,
		38905	=>	14581,
		38906	=>	14579,
		38907	=>	14576,
		38908	=>	14573,
		38909	=>	14571,
		38910	=>	14568,
		38911	=>	14565,
		38912	=>	14563,
		38913	=>	14560,
		38914	=>	14558,
		38915	=>	14555,
		38916	=>	14552,
		38917	=>	14550,
		38918	=>	14547,
		38919	=>	14545,
		38920	=>	14542,
		38921	=>	14539,
		38922	=>	14537,
		38923	=>	14534,
		38924	=>	14532,
		38925	=>	14529,
		38926	=>	14526,
		38927	=>	14524,
		38928	=>	14521,
		38929	=>	14518,
		38930	=>	14516,
		38931	=>	14513,
		38932	=>	14511,
		38933	=>	14508,
		38934	=>	14505,
		38935	=>	14503,
		38936	=>	14500,
		38937	=>	14498,
		38938	=>	14495,
		38939	=>	14492,
		38940	=>	14490,
		38941	=>	14487,
		38942	=>	14485,
		38943	=>	14482,
		38944	=>	14479,
		38945	=>	14477,
		38946	=>	14474,
		38947	=>	14472,
		38948	=>	14469,
		38949	=>	14466,
		38950	=>	14464,
		38951	=>	14461,
		38952	=>	14459,
		38953	=>	14456,
		38954	=>	14453,
		38955	=>	14451,
		38956	=>	14448,
		38957	=>	14445,
		38958	=>	14443,
		38959	=>	14440,
		38960	=>	14438,
		38961	=>	14435,
		38962	=>	14432,
		38963	=>	14430,
		38964	=>	14427,
		38965	=>	14425,
		38966	=>	14422,
		38967	=>	14419,
		38968	=>	14417,
		38969	=>	14414,
		38970	=>	14412,
		38971	=>	14409,
		38972	=>	14406,
		38973	=>	14404,
		38974	=>	14401,
		38975	=>	14399,
		38976	=>	14396,
		38977	=>	14393,
		38978	=>	14391,
		38979	=>	14388,
		38980	=>	14386,
		38981	=>	14383,
		38982	=>	14380,
		38983	=>	14378,
		38984	=>	14375,
		38985	=>	14373,
		38986	=>	14370,
		38987	=>	14367,
		38988	=>	14365,
		38989	=>	14362,
		38990	=>	14360,
		38991	=>	14357,
		38992	=>	14354,
		38993	=>	14352,
		38994	=>	14349,
		38995	=>	14347,
		38996	=>	14344,
		38997	=>	14341,
		38998	=>	14339,
		38999	=>	14336,
		39000	=>	14334,
		39001	=>	14331,
		39002	=>	14328,
		39003	=>	14326,
		39004	=>	14323,
		39005	=>	14321,
		39006	=>	14318,
		39007	=>	14315,
		39008	=>	14313,
		39009	=>	14310,
		39010	=>	14308,
		39011	=>	14305,
		39012	=>	14302,
		39013	=>	14300,
		39014	=>	14297,
		39015	=>	14295,
		39016	=>	14292,
		39017	=>	14290,
		39018	=>	14287,
		39019	=>	14284,
		39020	=>	14282,
		39021	=>	14279,
		39022	=>	14277,
		39023	=>	14274,
		39024	=>	14271,
		39025	=>	14269,
		39026	=>	14266,
		39027	=>	14264,
		39028	=>	14261,
		39029	=>	14258,
		39030	=>	14256,
		39031	=>	14253,
		39032	=>	14251,
		39033	=>	14248,
		39034	=>	14245,
		39035	=>	14243,
		39036	=>	14240,
		39037	=>	14238,
		39038	=>	14235,
		39039	=>	14232,
		39040	=>	14230,
		39041	=>	14227,
		39042	=>	14225,
		39043	=>	14222,
		39044	=>	14220,
		39045	=>	14217,
		39046	=>	14214,
		39047	=>	14212,
		39048	=>	14209,
		39049	=>	14207,
		39050	=>	14204,
		39051	=>	14201,
		39052	=>	14199,
		39053	=>	14196,
		39054	=>	14194,
		39055	=>	14191,
		39056	=>	14188,
		39057	=>	14186,
		39058	=>	14183,
		39059	=>	14181,
		39060	=>	14178,
		39061	=>	14176,
		39062	=>	14173,
		39063	=>	14170,
		39064	=>	14168,
		39065	=>	14165,
		39066	=>	14163,
		39067	=>	14160,
		39068	=>	14157,
		39069	=>	14155,
		39070	=>	14152,
		39071	=>	14150,
		39072	=>	14147,
		39073	=>	14144,
		39074	=>	14142,
		39075	=>	14139,
		39076	=>	14137,
		39077	=>	14134,
		39078	=>	14132,
		39079	=>	14129,
		39080	=>	14126,
		39081	=>	14124,
		39082	=>	14121,
		39083	=>	14119,
		39084	=>	14116,
		39085	=>	14113,
		39086	=>	14111,
		39087	=>	14108,
		39088	=>	14106,
		39089	=>	14103,
		39090	=>	14101,
		39091	=>	14098,
		39092	=>	14095,
		39093	=>	14093,
		39094	=>	14090,
		39095	=>	14088,
		39096	=>	14085,
		39097	=>	14083,
		39098	=>	14080,
		39099	=>	14077,
		39100	=>	14075,
		39101	=>	14072,
		39102	=>	14070,
		39103	=>	14067,
		39104	=>	14064,
		39105	=>	14062,
		39106	=>	14059,
		39107	=>	14057,
		39108	=>	14054,
		39109	=>	14052,
		39110	=>	14049,
		39111	=>	14046,
		39112	=>	14044,
		39113	=>	14041,
		39114	=>	14039,
		39115	=>	14036,
		39116	=>	14033,
		39117	=>	14031,
		39118	=>	14028,
		39119	=>	14026,
		39120	=>	14023,
		39121	=>	14021,
		39122	=>	14018,
		39123	=>	14015,
		39124	=>	14013,
		39125	=>	14010,
		39126	=>	14008,
		39127	=>	14005,
		39128	=>	14003,
		39129	=>	14000,
		39130	=>	13997,
		39131	=>	13995,
		39132	=>	13992,
		39133	=>	13990,
		39134	=>	13987,
		39135	=>	13985,
		39136	=>	13982,
		39137	=>	13979,
		39138	=>	13977,
		39139	=>	13974,
		39140	=>	13972,
		39141	=>	13969,
		39142	=>	13967,
		39143	=>	13964,
		39144	=>	13961,
		39145	=>	13959,
		39146	=>	13956,
		39147	=>	13954,
		39148	=>	13951,
		39149	=>	13949,
		39150	=>	13946,
		39151	=>	13943,
		39152	=>	13941,
		39153	=>	13938,
		39154	=>	13936,
		39155	=>	13933,
		39156	=>	13931,
		39157	=>	13928,
		39158	=>	13925,
		39159	=>	13923,
		39160	=>	13920,
		39161	=>	13918,
		39162	=>	13915,
		39163	=>	13913,
		39164	=>	13910,
		39165	=>	13907,
		39166	=>	13905,
		39167	=>	13902,
		39168	=>	13900,
		39169	=>	13897,
		39170	=>	13895,
		39171	=>	13892,
		39172	=>	13889,
		39173	=>	13887,
		39174	=>	13884,
		39175	=>	13882,
		39176	=>	13879,
		39177	=>	13877,
		39178	=>	13874,
		39179	=>	13871,
		39180	=>	13869,
		39181	=>	13866,
		39182	=>	13864,
		39183	=>	13861,
		39184	=>	13859,
		39185	=>	13856,
		39186	=>	13854,
		39187	=>	13851,
		39188	=>	13848,
		39189	=>	13846,
		39190	=>	13843,
		39191	=>	13841,
		39192	=>	13838,
		39193	=>	13836,
		39194	=>	13833,
		39195	=>	13830,
		39196	=>	13828,
		39197	=>	13825,
		39198	=>	13823,
		39199	=>	13820,
		39200	=>	13818,
		39201	=>	13815,
		39202	=>	13812,
		39203	=>	13810,
		39204	=>	13807,
		39205	=>	13805,
		39206	=>	13802,
		39207	=>	13800,
		39208	=>	13797,
		39209	=>	13795,
		39210	=>	13792,
		39211	=>	13789,
		39212	=>	13787,
		39213	=>	13784,
		39214	=>	13782,
		39215	=>	13779,
		39216	=>	13777,
		39217	=>	13774,
		39218	=>	13771,
		39219	=>	13769,
		39220	=>	13766,
		39221	=>	13764,
		39222	=>	13761,
		39223	=>	13759,
		39224	=>	13756,
		39225	=>	13754,
		39226	=>	13751,
		39227	=>	13748,
		39228	=>	13746,
		39229	=>	13743,
		39230	=>	13741,
		39231	=>	13738,
		39232	=>	13736,
		39233	=>	13733,
		39234	=>	13731,
		39235	=>	13728,
		39236	=>	13725,
		39237	=>	13723,
		39238	=>	13720,
		39239	=>	13718,
		39240	=>	13715,
		39241	=>	13713,
		39242	=>	13710,
		39243	=>	13708,
		39244	=>	13705,
		39245	=>	13702,
		39246	=>	13700,
		39247	=>	13697,
		39248	=>	13695,
		39249	=>	13692,
		39250	=>	13690,
		39251	=>	13687,
		39252	=>	13685,
		39253	=>	13682,
		39254	=>	13679,
		39255	=>	13677,
		39256	=>	13674,
		39257	=>	13672,
		39258	=>	13669,
		39259	=>	13667,
		39260	=>	13664,
		39261	=>	13662,
		39262	=>	13659,
		39263	=>	13656,
		39264	=>	13654,
		39265	=>	13651,
		39266	=>	13649,
		39267	=>	13646,
		39268	=>	13644,
		39269	=>	13641,
		39270	=>	13639,
		39271	=>	13636,
		39272	=>	13634,
		39273	=>	13631,
		39274	=>	13628,
		39275	=>	13626,
		39276	=>	13623,
		39277	=>	13621,
		39278	=>	13618,
		39279	=>	13616,
		39280	=>	13613,
		39281	=>	13611,
		39282	=>	13608,
		39283	=>	13605,
		39284	=>	13603,
		39285	=>	13600,
		39286	=>	13598,
		39287	=>	13595,
		39288	=>	13593,
		39289	=>	13590,
		39290	=>	13588,
		39291	=>	13585,
		39292	=>	13583,
		39293	=>	13580,
		39294	=>	13577,
		39295	=>	13575,
		39296	=>	13572,
		39297	=>	13570,
		39298	=>	13567,
		39299	=>	13565,
		39300	=>	13562,
		39301	=>	13560,
		39302	=>	13557,
		39303	=>	13555,
		39304	=>	13552,
		39305	=>	13549,
		39306	=>	13547,
		39307	=>	13544,
		39308	=>	13542,
		39309	=>	13539,
		39310	=>	13537,
		39311	=>	13534,
		39312	=>	13532,
		39313	=>	13529,
		39314	=>	13527,
		39315	=>	13524,
		39316	=>	13521,
		39317	=>	13519,
		39318	=>	13516,
		39319	=>	13514,
		39320	=>	13511,
		39321	=>	13509,
		39322	=>	13506,
		39323	=>	13504,
		39324	=>	13501,
		39325	=>	13499,
		39326	=>	13496,
		39327	=>	13494,
		39328	=>	13491,
		39329	=>	13488,
		39330	=>	13486,
		39331	=>	13483,
		39332	=>	13481,
		39333	=>	13478,
		39334	=>	13476,
		39335	=>	13473,
		39336	=>	13471,
		39337	=>	13468,
		39338	=>	13466,
		39339	=>	13463,
		39340	=>	13461,
		39341	=>	13458,
		39342	=>	13455,
		39343	=>	13453,
		39344	=>	13450,
		39345	=>	13448,
		39346	=>	13445,
		39347	=>	13443,
		39348	=>	13440,
		39349	=>	13438,
		39350	=>	13435,
		39351	=>	13433,
		39352	=>	13430,
		39353	=>	13428,
		39354	=>	13425,
		39355	=>	13422,
		39356	=>	13420,
		39357	=>	13417,
		39358	=>	13415,
		39359	=>	13412,
		39360	=>	13410,
		39361	=>	13407,
		39362	=>	13405,
		39363	=>	13402,
		39364	=>	13400,
		39365	=>	13397,
		39366	=>	13395,
		39367	=>	13392,
		39368	=>	13390,
		39369	=>	13387,
		39370	=>	13384,
		39371	=>	13382,
		39372	=>	13379,
		39373	=>	13377,
		39374	=>	13374,
		39375	=>	13372,
		39376	=>	13369,
		39377	=>	13367,
		39378	=>	13364,
		39379	=>	13362,
		39380	=>	13359,
		39381	=>	13357,
		39382	=>	13354,
		39383	=>	13352,
		39384	=>	13349,
		39385	=>	13346,
		39386	=>	13344,
		39387	=>	13341,
		39388	=>	13339,
		39389	=>	13336,
		39390	=>	13334,
		39391	=>	13331,
		39392	=>	13329,
		39393	=>	13326,
		39394	=>	13324,
		39395	=>	13321,
		39396	=>	13319,
		39397	=>	13316,
		39398	=>	13314,
		39399	=>	13311,
		39400	=>	13309,
		39401	=>	13306,
		39402	=>	13303,
		39403	=>	13301,
		39404	=>	13298,
		39405	=>	13296,
		39406	=>	13293,
		39407	=>	13291,
		39408	=>	13288,
		39409	=>	13286,
		39410	=>	13283,
		39411	=>	13281,
		39412	=>	13278,
		39413	=>	13276,
		39414	=>	13273,
		39415	=>	13271,
		39416	=>	13268,
		39417	=>	13266,
		39418	=>	13263,
		39419	=>	13261,
		39420	=>	13258,
		39421	=>	13255,
		39422	=>	13253,
		39423	=>	13250,
		39424	=>	13248,
		39425	=>	13245,
		39426	=>	13243,
		39427	=>	13240,
		39428	=>	13238,
		39429	=>	13235,
		39430	=>	13233,
		39431	=>	13230,
		39432	=>	13228,
		39433	=>	13225,
		39434	=>	13223,
		39435	=>	13220,
		39436	=>	13218,
		39437	=>	13215,
		39438	=>	13213,
		39439	=>	13210,
		39440	=>	13208,
		39441	=>	13205,
		39442	=>	13203,
		39443	=>	13200,
		39444	=>	13197,
		39445	=>	13195,
		39446	=>	13192,
		39447	=>	13190,
		39448	=>	13187,
		39449	=>	13185,
		39450	=>	13182,
		39451	=>	13180,
		39452	=>	13177,
		39453	=>	13175,
		39454	=>	13172,
		39455	=>	13170,
		39456	=>	13167,
		39457	=>	13165,
		39458	=>	13162,
		39459	=>	13160,
		39460	=>	13157,
		39461	=>	13155,
		39462	=>	13152,
		39463	=>	13150,
		39464	=>	13147,
		39465	=>	13145,
		39466	=>	13142,
		39467	=>	13140,
		39468	=>	13137,
		39469	=>	13135,
		39470	=>	13132,
		39471	=>	13130,
		39472	=>	13127,
		39473	=>	13124,
		39474	=>	13122,
		39475	=>	13119,
		39476	=>	13117,
		39477	=>	13114,
		39478	=>	13112,
		39479	=>	13109,
		39480	=>	13107,
		39481	=>	13104,
		39482	=>	13102,
		39483	=>	13099,
		39484	=>	13097,
		39485	=>	13094,
		39486	=>	13092,
		39487	=>	13089,
		39488	=>	13087,
		39489	=>	13084,
		39490	=>	13082,
		39491	=>	13079,
		39492	=>	13077,
		39493	=>	13074,
		39494	=>	13072,
		39495	=>	13069,
		39496	=>	13067,
		39497	=>	13064,
		39498	=>	13062,
		39499	=>	13059,
		39500	=>	13057,
		39501	=>	13054,
		39502	=>	13052,
		39503	=>	13049,
		39504	=>	13047,
		39505	=>	13044,
		39506	=>	13042,
		39507	=>	13039,
		39508	=>	13037,
		39509	=>	13034,
		39510	=>	13032,
		39511	=>	13029,
		39512	=>	13027,
		39513	=>	13024,
		39514	=>	13022,
		39515	=>	13019,
		39516	=>	13017,
		39517	=>	13014,
		39518	=>	13012,
		39519	=>	13009,
		39520	=>	13007,
		39521	=>	13004,
		39522	=>	13002,
		39523	=>	12999,
		39524	=>	12996,
		39525	=>	12994,
		39526	=>	12991,
		39527	=>	12989,
		39528	=>	12986,
		39529	=>	12984,
		39530	=>	12981,
		39531	=>	12979,
		39532	=>	12976,
		39533	=>	12974,
		39534	=>	12971,
		39535	=>	12969,
		39536	=>	12966,
		39537	=>	12964,
		39538	=>	12961,
		39539	=>	12959,
		39540	=>	12956,
		39541	=>	12954,
		39542	=>	12951,
		39543	=>	12949,
		39544	=>	12946,
		39545	=>	12944,
		39546	=>	12941,
		39547	=>	12939,
		39548	=>	12936,
		39549	=>	12934,
		39550	=>	12931,
		39551	=>	12929,
		39552	=>	12926,
		39553	=>	12924,
		39554	=>	12921,
		39555	=>	12919,
		39556	=>	12916,
		39557	=>	12914,
		39558	=>	12911,
		39559	=>	12909,
		39560	=>	12906,
		39561	=>	12904,
		39562	=>	12901,
		39563	=>	12899,
		39564	=>	12896,
		39565	=>	12894,
		39566	=>	12891,
		39567	=>	12889,
		39568	=>	12886,
		39569	=>	12884,
		39570	=>	12881,
		39571	=>	12879,
		39572	=>	12876,
		39573	=>	12874,
		39574	=>	12871,
		39575	=>	12869,
		39576	=>	12866,
		39577	=>	12864,
		39578	=>	12861,
		39579	=>	12859,
		39580	=>	12856,
		39581	=>	12854,
		39582	=>	12851,
		39583	=>	12849,
		39584	=>	12847,
		39585	=>	12844,
		39586	=>	12842,
		39587	=>	12839,
		39588	=>	12837,
		39589	=>	12834,
		39590	=>	12832,
		39591	=>	12829,
		39592	=>	12827,
		39593	=>	12824,
		39594	=>	12822,
		39595	=>	12819,
		39596	=>	12817,
		39597	=>	12814,
		39598	=>	12812,
		39599	=>	12809,
		39600	=>	12807,
		39601	=>	12804,
		39602	=>	12802,
		39603	=>	12799,
		39604	=>	12797,
		39605	=>	12794,
		39606	=>	12792,
		39607	=>	12789,
		39608	=>	12787,
		39609	=>	12784,
		39610	=>	12782,
		39611	=>	12779,
		39612	=>	12777,
		39613	=>	12774,
		39614	=>	12772,
		39615	=>	12769,
		39616	=>	12767,
		39617	=>	12764,
		39618	=>	12762,
		39619	=>	12759,
		39620	=>	12757,
		39621	=>	12754,
		39622	=>	12752,
		39623	=>	12749,
		39624	=>	12747,
		39625	=>	12744,
		39626	=>	12742,
		39627	=>	12739,
		39628	=>	12737,
		39629	=>	12734,
		39630	=>	12732,
		39631	=>	12729,
		39632	=>	12727,
		39633	=>	12725,
		39634	=>	12722,
		39635	=>	12720,
		39636	=>	12717,
		39637	=>	12715,
		39638	=>	12712,
		39639	=>	12710,
		39640	=>	12707,
		39641	=>	12705,
		39642	=>	12702,
		39643	=>	12700,
		39644	=>	12697,
		39645	=>	12695,
		39646	=>	12692,
		39647	=>	12690,
		39648	=>	12687,
		39649	=>	12685,
		39650	=>	12682,
		39651	=>	12680,
		39652	=>	12677,
		39653	=>	12675,
		39654	=>	12672,
		39655	=>	12670,
		39656	=>	12667,
		39657	=>	12665,
		39658	=>	12662,
		39659	=>	12660,
		39660	=>	12657,
		39661	=>	12655,
		39662	=>	12653,
		39663	=>	12650,
		39664	=>	12648,
		39665	=>	12645,
		39666	=>	12643,
		39667	=>	12640,
		39668	=>	12638,
		39669	=>	12635,
		39670	=>	12633,
		39671	=>	12630,
		39672	=>	12628,
		39673	=>	12625,
		39674	=>	12623,
		39675	=>	12620,
		39676	=>	12618,
		39677	=>	12615,
		39678	=>	12613,
		39679	=>	12610,
		39680	=>	12608,
		39681	=>	12605,
		39682	=>	12603,
		39683	=>	12600,
		39684	=>	12598,
		39685	=>	12596,
		39686	=>	12593,
		39687	=>	12591,
		39688	=>	12588,
		39689	=>	12586,
		39690	=>	12583,
		39691	=>	12581,
		39692	=>	12578,
		39693	=>	12576,
		39694	=>	12573,
		39695	=>	12571,
		39696	=>	12568,
		39697	=>	12566,
		39698	=>	12563,
		39699	=>	12561,
		39700	=>	12558,
		39701	=>	12556,
		39702	=>	12553,
		39703	=>	12551,
		39704	=>	12549,
		39705	=>	12546,
		39706	=>	12544,
		39707	=>	12541,
		39708	=>	12539,
		39709	=>	12536,
		39710	=>	12534,
		39711	=>	12531,
		39712	=>	12529,
		39713	=>	12526,
		39714	=>	12524,
		39715	=>	12521,
		39716	=>	12519,
		39717	=>	12516,
		39718	=>	12514,
		39719	=>	12511,
		39720	=>	12509,
		39721	=>	12507,
		39722	=>	12504,
		39723	=>	12502,
		39724	=>	12499,
		39725	=>	12497,
		39726	=>	12494,
		39727	=>	12492,
		39728	=>	12489,
		39729	=>	12487,
		39730	=>	12484,
		39731	=>	12482,
		39732	=>	12479,
		39733	=>	12477,
		39734	=>	12474,
		39735	=>	12472,
		39736	=>	12469,
		39737	=>	12467,
		39738	=>	12465,
		39739	=>	12462,
		39740	=>	12460,
		39741	=>	12457,
		39742	=>	12455,
		39743	=>	12452,
		39744	=>	12450,
		39745	=>	12447,
		39746	=>	12445,
		39747	=>	12442,
		39748	=>	12440,
		39749	=>	12437,
		39750	=>	12435,
		39751	=>	12433,
		39752	=>	12430,
		39753	=>	12428,
		39754	=>	12425,
		39755	=>	12423,
		39756	=>	12420,
		39757	=>	12418,
		39758	=>	12415,
		39759	=>	12413,
		39760	=>	12410,
		39761	=>	12408,
		39762	=>	12405,
		39763	=>	12403,
		39764	=>	12401,
		39765	=>	12398,
		39766	=>	12396,
		39767	=>	12393,
		39768	=>	12391,
		39769	=>	12388,
		39770	=>	12386,
		39771	=>	12383,
		39772	=>	12381,
		39773	=>	12378,
		39774	=>	12376,
		39775	=>	12373,
		39776	=>	12371,
		39777	=>	12369,
		39778	=>	12366,
		39779	=>	12364,
		39780	=>	12361,
		39781	=>	12359,
		39782	=>	12356,
		39783	=>	12354,
		39784	=>	12351,
		39785	=>	12349,
		39786	=>	12346,
		39787	=>	12344,
		39788	=>	12342,
		39789	=>	12339,
		39790	=>	12337,
		39791	=>	12334,
		39792	=>	12332,
		39793	=>	12329,
		39794	=>	12327,
		39795	=>	12324,
		39796	=>	12322,
		39797	=>	12319,
		39798	=>	12317,
		39799	=>	12314,
		39800	=>	12312,
		39801	=>	12310,
		39802	=>	12307,
		39803	=>	12305,
		39804	=>	12302,
		39805	=>	12300,
		39806	=>	12297,
		39807	=>	12295,
		39808	=>	12292,
		39809	=>	12290,
		39810	=>	12288,
		39811	=>	12285,
		39812	=>	12283,
		39813	=>	12280,
		39814	=>	12278,
		39815	=>	12275,
		39816	=>	12273,
		39817	=>	12270,
		39818	=>	12268,
		39819	=>	12265,
		39820	=>	12263,
		39821	=>	12261,
		39822	=>	12258,
		39823	=>	12256,
		39824	=>	12253,
		39825	=>	12251,
		39826	=>	12248,
		39827	=>	12246,
		39828	=>	12243,
		39829	=>	12241,
		39830	=>	12239,
		39831	=>	12236,
		39832	=>	12234,
		39833	=>	12231,
		39834	=>	12229,
		39835	=>	12226,
		39836	=>	12224,
		39837	=>	12221,
		39838	=>	12219,
		39839	=>	12216,
		39840	=>	12214,
		39841	=>	12212,
		39842	=>	12209,
		39843	=>	12207,
		39844	=>	12204,
		39845	=>	12202,
		39846	=>	12199,
		39847	=>	12197,
		39848	=>	12194,
		39849	=>	12192,
		39850	=>	12190,
		39851	=>	12187,
		39852	=>	12185,
		39853	=>	12182,
		39854	=>	12180,
		39855	=>	12177,
		39856	=>	12175,
		39857	=>	12172,
		39858	=>	12170,
		39859	=>	12168,
		39860	=>	12165,
		39861	=>	12163,
		39862	=>	12160,
		39863	=>	12158,
		39864	=>	12155,
		39865	=>	12153,
		39866	=>	12150,
		39867	=>	12148,
		39868	=>	12146,
		39869	=>	12143,
		39870	=>	12141,
		39871	=>	12138,
		39872	=>	12136,
		39873	=>	12133,
		39874	=>	12131,
		39875	=>	12129,
		39876	=>	12126,
		39877	=>	12124,
		39878	=>	12121,
		39879	=>	12119,
		39880	=>	12116,
		39881	=>	12114,
		39882	=>	12111,
		39883	=>	12109,
		39884	=>	12107,
		39885	=>	12104,
		39886	=>	12102,
		39887	=>	12099,
		39888	=>	12097,
		39889	=>	12094,
		39890	=>	12092,
		39891	=>	12089,
		39892	=>	12087,
		39893	=>	12085,
		39894	=>	12082,
		39895	=>	12080,
		39896	=>	12077,
		39897	=>	12075,
		39898	=>	12072,
		39899	=>	12070,
		39900	=>	12068,
		39901	=>	12065,
		39902	=>	12063,
		39903	=>	12060,
		39904	=>	12058,
		39905	=>	12055,
		39906	=>	12053,
		39907	=>	12051,
		39908	=>	12048,
		39909	=>	12046,
		39910	=>	12043,
		39911	=>	12041,
		39912	=>	12038,
		39913	=>	12036,
		39914	=>	12033,
		39915	=>	12031,
		39916	=>	12029,
		39917	=>	12026,
		39918	=>	12024,
		39919	=>	12021,
		39920	=>	12019,
		39921	=>	12016,
		39922	=>	12014,
		39923	=>	12012,
		39924	=>	12009,
		39925	=>	12007,
		39926	=>	12004,
		39927	=>	12002,
		39928	=>	11999,
		39929	=>	11997,
		39930	=>	11995,
		39931	=>	11992,
		39932	=>	11990,
		39933	=>	11987,
		39934	=>	11985,
		39935	=>	11982,
		39936	=>	11980,
		39937	=>	11978,
		39938	=>	11975,
		39939	=>	11973,
		39940	=>	11970,
		39941	=>	11968,
		39942	=>	11965,
		39943	=>	11963,
		39944	=>	11961,
		39945	=>	11958,
		39946	=>	11956,
		39947	=>	11953,
		39948	=>	11951,
		39949	=>	11948,
		39950	=>	11946,
		39951	=>	11944,
		39952	=>	11941,
		39953	=>	11939,
		39954	=>	11936,
		39955	=>	11934,
		39956	=>	11931,
		39957	=>	11929,
		39958	=>	11927,
		39959	=>	11924,
		39960	=>	11922,
		39961	=>	11919,
		39962	=>	11917,
		39963	=>	11915,
		39964	=>	11912,
		39965	=>	11910,
		39966	=>	11907,
		39967	=>	11905,
		39968	=>	11902,
		39969	=>	11900,
		39970	=>	11898,
		39971	=>	11895,
		39972	=>	11893,
		39973	=>	11890,
		39974	=>	11888,
		39975	=>	11885,
		39976	=>	11883,
		39977	=>	11881,
		39978	=>	11878,
		39979	=>	11876,
		39980	=>	11873,
		39981	=>	11871,
		39982	=>	11869,
		39983	=>	11866,
		39984	=>	11864,
		39985	=>	11861,
		39986	=>	11859,
		39987	=>	11856,
		39988	=>	11854,
		39989	=>	11852,
		39990	=>	11849,
		39991	=>	11847,
		39992	=>	11844,
		39993	=>	11842,
		39994	=>	11839,
		39995	=>	11837,
		39996	=>	11835,
		39997	=>	11832,
		39998	=>	11830,
		39999	=>	11827,
		40000	=>	11825,
		40001	=>	11823,
		40002	=>	11820,
		40003	=>	11818,
		40004	=>	11815,
		40005	=>	11813,
		40006	=>	11810,
		40007	=>	11808,
		40008	=>	11806,
		40009	=>	11803,
		40010	=>	11801,
		40011	=>	11798,
		40012	=>	11796,
		40013	=>	11794,
		40014	=>	11791,
		40015	=>	11789,
		40016	=>	11786,
		40017	=>	11784,
		40018	=>	11782,
		40019	=>	11779,
		40020	=>	11777,
		40021	=>	11774,
		40022	=>	11772,
		40023	=>	11769,
		40024	=>	11767,
		40025	=>	11765,
		40026	=>	11762,
		40027	=>	11760,
		40028	=>	11757,
		40029	=>	11755,
		40030	=>	11753,
		40031	=>	11750,
		40032	=>	11748,
		40033	=>	11745,
		40034	=>	11743,
		40035	=>	11741,
		40036	=>	11738,
		40037	=>	11736,
		40038	=>	11733,
		40039	=>	11731,
		40040	=>	11728,
		40041	=>	11726,
		40042	=>	11724,
		40043	=>	11721,
		40044	=>	11719,
		40045	=>	11716,
		40046	=>	11714,
		40047	=>	11712,
		40048	=>	11709,
		40049	=>	11707,
		40050	=>	11704,
		40051	=>	11702,
		40052	=>	11700,
		40053	=>	11697,
		40054	=>	11695,
		40055	=>	11692,
		40056	=>	11690,
		40057	=>	11688,
		40058	=>	11685,
		40059	=>	11683,
		40060	=>	11680,
		40061	=>	11678,
		40062	=>	11676,
		40063	=>	11673,
		40064	=>	11671,
		40065	=>	11668,
		40066	=>	11666,
		40067	=>	11664,
		40068	=>	11661,
		40069	=>	11659,
		40070	=>	11656,
		40071	=>	11654,
		40072	=>	11652,
		40073	=>	11649,
		40074	=>	11647,
		40075	=>	11644,
		40076	=>	11642,
		40077	=>	11640,
		40078	=>	11637,
		40079	=>	11635,
		40080	=>	11632,
		40081	=>	11630,
		40082	=>	11628,
		40083	=>	11625,
		40084	=>	11623,
		40085	=>	11620,
		40086	=>	11618,
		40087	=>	11616,
		40088	=>	11613,
		40089	=>	11611,
		40090	=>	11608,
		40091	=>	11606,
		40092	=>	11604,
		40093	=>	11601,
		40094	=>	11599,
		40095	=>	11596,
		40096	=>	11594,
		40097	=>	11592,
		40098	=>	11589,
		40099	=>	11587,
		40100	=>	11584,
		40101	=>	11582,
		40102	=>	11580,
		40103	=>	11577,
		40104	=>	11575,
		40105	=>	11572,
		40106	=>	11570,
		40107	=>	11568,
		40108	=>	11565,
		40109	=>	11563,
		40110	=>	11560,
		40111	=>	11558,
		40112	=>	11556,
		40113	=>	11553,
		40114	=>	11551,
		40115	=>	11548,
		40116	=>	11546,
		40117	=>	11544,
		40118	=>	11541,
		40119	=>	11539,
		40120	=>	11536,
		40121	=>	11534,
		40122	=>	11532,
		40123	=>	11529,
		40124	=>	11527,
		40125	=>	11524,
		40126	=>	11522,
		40127	=>	11520,
		40128	=>	11517,
		40129	=>	11515,
		40130	=>	11513,
		40131	=>	11510,
		40132	=>	11508,
		40133	=>	11505,
		40134	=>	11503,
		40135	=>	11501,
		40136	=>	11498,
		40137	=>	11496,
		40138	=>	11493,
		40139	=>	11491,
		40140	=>	11489,
		40141	=>	11486,
		40142	=>	11484,
		40143	=>	11481,
		40144	=>	11479,
		40145	=>	11477,
		40146	=>	11474,
		40147	=>	11472,
		40148	=>	11470,
		40149	=>	11467,
		40150	=>	11465,
		40151	=>	11462,
		40152	=>	11460,
		40153	=>	11458,
		40154	=>	11455,
		40155	=>	11453,
		40156	=>	11450,
		40157	=>	11448,
		40158	=>	11446,
		40159	=>	11443,
		40160	=>	11441,
		40161	=>	11438,
		40162	=>	11436,
		40163	=>	11434,
		40164	=>	11431,
		40165	=>	11429,
		40166	=>	11427,
		40167	=>	11424,
		40168	=>	11422,
		40169	=>	11419,
		40170	=>	11417,
		40171	=>	11415,
		40172	=>	11412,
		40173	=>	11410,
		40174	=>	11408,
		40175	=>	11405,
		40176	=>	11403,
		40177	=>	11400,
		40178	=>	11398,
		40179	=>	11396,
		40180	=>	11393,
		40181	=>	11391,
		40182	=>	11388,
		40183	=>	11386,
		40184	=>	11384,
		40185	=>	11381,
		40186	=>	11379,
		40187	=>	11377,
		40188	=>	11374,
		40189	=>	11372,
		40190	=>	11369,
		40191	=>	11367,
		40192	=>	11365,
		40193	=>	11362,
		40194	=>	11360,
		40195	=>	11358,
		40196	=>	11355,
		40197	=>	11353,
		40198	=>	11350,
		40199	=>	11348,
		40200	=>	11346,
		40201	=>	11343,
		40202	=>	11341,
		40203	=>	11339,
		40204	=>	11336,
		40205	=>	11334,
		40206	=>	11331,
		40207	=>	11329,
		40208	=>	11327,
		40209	=>	11324,
		40210	=>	11322,
		40211	=>	11319,
		40212	=>	11317,
		40213	=>	11315,
		40214	=>	11312,
		40215	=>	11310,
		40216	=>	11308,
		40217	=>	11305,
		40218	=>	11303,
		40219	=>	11301,
		40220	=>	11298,
		40221	=>	11296,
		40222	=>	11293,
		40223	=>	11291,
		40224	=>	11289,
		40225	=>	11286,
		40226	=>	11284,
		40227	=>	11282,
		40228	=>	11279,
		40229	=>	11277,
		40230	=>	11274,
		40231	=>	11272,
		40232	=>	11270,
		40233	=>	11267,
		40234	=>	11265,
		40235	=>	11263,
		40236	=>	11260,
		40237	=>	11258,
		40238	=>	11255,
		40239	=>	11253,
		40240	=>	11251,
		40241	=>	11248,
		40242	=>	11246,
		40243	=>	11244,
		40244	=>	11241,
		40245	=>	11239,
		40246	=>	11236,
		40247	=>	11234,
		40248	=>	11232,
		40249	=>	11229,
		40250	=>	11227,
		40251	=>	11225,
		40252	=>	11222,
		40253	=>	11220,
		40254	=>	11218,
		40255	=>	11215,
		40256	=>	11213,
		40257	=>	11210,
		40258	=>	11208,
		40259	=>	11206,
		40260	=>	11203,
		40261	=>	11201,
		40262	=>	11199,
		40263	=>	11196,
		40264	=>	11194,
		40265	=>	11192,
		40266	=>	11189,
		40267	=>	11187,
		40268	=>	11184,
		40269	=>	11182,
		40270	=>	11180,
		40271	=>	11177,
		40272	=>	11175,
		40273	=>	11173,
		40274	=>	11170,
		40275	=>	11168,
		40276	=>	11166,
		40277	=>	11163,
		40278	=>	11161,
		40279	=>	11158,
		40280	=>	11156,
		40281	=>	11154,
		40282	=>	11151,
		40283	=>	11149,
		40284	=>	11147,
		40285	=>	11144,
		40286	=>	11142,
		40287	=>	11140,
		40288	=>	11137,
		40289	=>	11135,
		40290	=>	11132,
		40291	=>	11130,
		40292	=>	11128,
		40293	=>	11125,
		40294	=>	11123,
		40295	=>	11121,
		40296	=>	11118,
		40297	=>	11116,
		40298	=>	11114,
		40299	=>	11111,
		40300	=>	11109,
		40301	=>	11107,
		40302	=>	11104,
		40303	=>	11102,
		40304	=>	11099,
		40305	=>	11097,
		40306	=>	11095,
		40307	=>	11092,
		40308	=>	11090,
		40309	=>	11088,
		40310	=>	11085,
		40311	=>	11083,
		40312	=>	11081,
		40313	=>	11078,
		40314	=>	11076,
		40315	=>	11074,
		40316	=>	11071,
		40317	=>	11069,
		40318	=>	11066,
		40319	=>	11064,
		40320	=>	11062,
		40321	=>	11059,
		40322	=>	11057,
		40323	=>	11055,
		40324	=>	11052,
		40325	=>	11050,
		40326	=>	11048,
		40327	=>	11045,
		40328	=>	11043,
		40329	=>	11041,
		40330	=>	11038,
		40331	=>	11036,
		40332	=>	11034,
		40333	=>	11031,
		40334	=>	11029,
		40335	=>	11027,
		40336	=>	11024,
		40337	=>	11022,
		40338	=>	11019,
		40339	=>	11017,
		40340	=>	11015,
		40341	=>	11012,
		40342	=>	11010,
		40343	=>	11008,
		40344	=>	11005,
		40345	=>	11003,
		40346	=>	11001,
		40347	=>	10998,
		40348	=>	10996,
		40349	=>	10994,
		40350	=>	10991,
		40351	=>	10989,
		40352	=>	10987,
		40353	=>	10984,
		40354	=>	10982,
		40355	=>	10980,
		40356	=>	10977,
		40357	=>	10975,
		40358	=>	10973,
		40359	=>	10970,
		40360	=>	10968,
		40361	=>	10965,
		40362	=>	10963,
		40363	=>	10961,
		40364	=>	10958,
		40365	=>	10956,
		40366	=>	10954,
		40367	=>	10951,
		40368	=>	10949,
		40369	=>	10947,
		40370	=>	10944,
		40371	=>	10942,
		40372	=>	10940,
		40373	=>	10937,
		40374	=>	10935,
		40375	=>	10933,
		40376	=>	10930,
		40377	=>	10928,
		40378	=>	10926,
		40379	=>	10923,
		40380	=>	10921,
		40381	=>	10919,
		40382	=>	10916,
		40383	=>	10914,
		40384	=>	10912,
		40385	=>	10909,
		40386	=>	10907,
		40387	=>	10905,
		40388	=>	10902,
		40389	=>	10900,
		40390	=>	10898,
		40391	=>	10895,
		40392	=>	10893,
		40393	=>	10891,
		40394	=>	10888,
		40395	=>	10886,
		40396	=>	10884,
		40397	=>	10881,
		40398	=>	10879,
		40399	=>	10876,
		40400	=>	10874,
		40401	=>	10872,
		40402	=>	10869,
		40403	=>	10867,
		40404	=>	10865,
		40405	=>	10862,
		40406	=>	10860,
		40407	=>	10858,
		40408	=>	10855,
		40409	=>	10853,
		40410	=>	10851,
		40411	=>	10848,
		40412	=>	10846,
		40413	=>	10844,
		40414	=>	10841,
		40415	=>	10839,
		40416	=>	10837,
		40417	=>	10834,
		40418	=>	10832,
		40419	=>	10830,
		40420	=>	10827,
		40421	=>	10825,
		40422	=>	10823,
		40423	=>	10820,
		40424	=>	10818,
		40425	=>	10816,
		40426	=>	10813,
		40427	=>	10811,
		40428	=>	10809,
		40429	=>	10806,
		40430	=>	10804,
		40431	=>	10802,
		40432	=>	10799,
		40433	=>	10797,
		40434	=>	10795,
		40435	=>	10792,
		40436	=>	10790,
		40437	=>	10788,
		40438	=>	10785,
		40439	=>	10783,
		40440	=>	10781,
		40441	=>	10778,
		40442	=>	10776,
		40443	=>	10774,
		40444	=>	10772,
		40445	=>	10769,
		40446	=>	10767,
		40447	=>	10765,
		40448	=>	10762,
		40449	=>	10760,
		40450	=>	10758,
		40451	=>	10755,
		40452	=>	10753,
		40453	=>	10751,
		40454	=>	10748,
		40455	=>	10746,
		40456	=>	10744,
		40457	=>	10741,
		40458	=>	10739,
		40459	=>	10737,
		40460	=>	10734,
		40461	=>	10732,
		40462	=>	10730,
		40463	=>	10727,
		40464	=>	10725,
		40465	=>	10723,
		40466	=>	10720,
		40467	=>	10718,
		40468	=>	10716,
		40469	=>	10713,
		40470	=>	10711,
		40471	=>	10709,
		40472	=>	10706,
		40473	=>	10704,
		40474	=>	10702,
		40475	=>	10699,
		40476	=>	10697,
		40477	=>	10695,
		40478	=>	10692,
		40479	=>	10690,
		40480	=>	10688,
		40481	=>	10685,
		40482	=>	10683,
		40483	=>	10681,
		40484	=>	10679,
		40485	=>	10676,
		40486	=>	10674,
		40487	=>	10672,
		40488	=>	10669,
		40489	=>	10667,
		40490	=>	10665,
		40491	=>	10662,
		40492	=>	10660,
		40493	=>	10658,
		40494	=>	10655,
		40495	=>	10653,
		40496	=>	10651,
		40497	=>	10648,
		40498	=>	10646,
		40499	=>	10644,
		40500	=>	10641,
		40501	=>	10639,
		40502	=>	10637,
		40503	=>	10634,
		40504	=>	10632,
		40505	=>	10630,
		40506	=>	10628,
		40507	=>	10625,
		40508	=>	10623,
		40509	=>	10621,
		40510	=>	10618,
		40511	=>	10616,
		40512	=>	10614,
		40513	=>	10611,
		40514	=>	10609,
		40515	=>	10607,
		40516	=>	10604,
		40517	=>	10602,
		40518	=>	10600,
		40519	=>	10597,
		40520	=>	10595,
		40521	=>	10593,
		40522	=>	10590,
		40523	=>	10588,
		40524	=>	10586,
		40525	=>	10584,
		40526	=>	10581,
		40527	=>	10579,
		40528	=>	10577,
		40529	=>	10574,
		40530	=>	10572,
		40531	=>	10570,
		40532	=>	10567,
		40533	=>	10565,
		40534	=>	10563,
		40535	=>	10560,
		40536	=>	10558,
		40537	=>	10556,
		40538	=>	10554,
		40539	=>	10551,
		40540	=>	10549,
		40541	=>	10547,
		40542	=>	10544,
		40543	=>	10542,
		40544	=>	10540,
		40545	=>	10537,
		40546	=>	10535,
		40547	=>	10533,
		40548	=>	10530,
		40549	=>	10528,
		40550	=>	10526,
		40551	=>	10524,
		40552	=>	10521,
		40553	=>	10519,
		40554	=>	10517,
		40555	=>	10514,
		40556	=>	10512,
		40557	=>	10510,
		40558	=>	10507,
		40559	=>	10505,
		40560	=>	10503,
		40561	=>	10500,
		40562	=>	10498,
		40563	=>	10496,
		40564	=>	10494,
		40565	=>	10491,
		40566	=>	10489,
		40567	=>	10487,
		40568	=>	10484,
		40569	=>	10482,
		40570	=>	10480,
		40571	=>	10477,
		40572	=>	10475,
		40573	=>	10473,
		40574	=>	10471,
		40575	=>	10468,
		40576	=>	10466,
		40577	=>	10464,
		40578	=>	10461,
		40579	=>	10459,
		40580	=>	10457,
		40581	=>	10454,
		40582	=>	10452,
		40583	=>	10450,
		40584	=>	10448,
		40585	=>	10445,
		40586	=>	10443,
		40587	=>	10441,
		40588	=>	10438,
		40589	=>	10436,
		40590	=>	10434,
		40591	=>	10431,
		40592	=>	10429,
		40593	=>	10427,
		40594	=>	10425,
		40595	=>	10422,
		40596	=>	10420,
		40597	=>	10418,
		40598	=>	10415,
		40599	=>	10413,
		40600	=>	10411,
		40601	=>	10408,
		40602	=>	10406,
		40603	=>	10404,
		40604	=>	10402,
		40605	=>	10399,
		40606	=>	10397,
		40607	=>	10395,
		40608	=>	10392,
		40609	=>	10390,
		40610	=>	10388,
		40611	=>	10385,
		40612	=>	10383,
		40613	=>	10381,
		40614	=>	10379,
		40615	=>	10376,
		40616	=>	10374,
		40617	=>	10372,
		40618	=>	10369,
		40619	=>	10367,
		40620	=>	10365,
		40621	=>	10363,
		40622	=>	10360,
		40623	=>	10358,
		40624	=>	10356,
		40625	=>	10353,
		40626	=>	10351,
		40627	=>	10349,
		40628	=>	10346,
		40629	=>	10344,
		40630	=>	10342,
		40631	=>	10340,
		40632	=>	10337,
		40633	=>	10335,
		40634	=>	10333,
		40635	=>	10330,
		40636	=>	10328,
		40637	=>	10326,
		40638	=>	10324,
		40639	=>	10321,
		40640	=>	10319,
		40641	=>	10317,
		40642	=>	10314,
		40643	=>	10312,
		40644	=>	10310,
		40645	=>	10308,
		40646	=>	10305,
		40647	=>	10303,
		40648	=>	10301,
		40649	=>	10298,
		40650	=>	10296,
		40651	=>	10294,
		40652	=>	10292,
		40653	=>	10289,
		40654	=>	10287,
		40655	=>	10285,
		40656	=>	10282,
		40657	=>	10280,
		40658	=>	10278,
		40659	=>	10276,
		40660	=>	10273,
		40661	=>	10271,
		40662	=>	10269,
		40663	=>	10266,
		40664	=>	10264,
		40665	=>	10262,
		40666	=>	10260,
		40667	=>	10257,
		40668	=>	10255,
		40669	=>	10253,
		40670	=>	10250,
		40671	=>	10248,
		40672	=>	10246,
		40673	=>	10244,
		40674	=>	10241,
		40675	=>	10239,
		40676	=>	10237,
		40677	=>	10234,
		40678	=>	10232,
		40679	=>	10230,
		40680	=>	10228,
		40681	=>	10225,
		40682	=>	10223,
		40683	=>	10221,
		40684	=>	10219,
		40685	=>	10216,
		40686	=>	10214,
		40687	=>	10212,
		40688	=>	10209,
		40689	=>	10207,
		40690	=>	10205,
		40691	=>	10203,
		40692	=>	10200,
		40693	=>	10198,
		40694	=>	10196,
		40695	=>	10193,
		40696	=>	10191,
		40697	=>	10189,
		40698	=>	10187,
		40699	=>	10184,
		40700	=>	10182,
		40701	=>	10180,
		40702	=>	10178,
		40703	=>	10175,
		40704	=>	10173,
		40705	=>	10171,
		40706	=>	10168,
		40707	=>	10166,
		40708	=>	10164,
		40709	=>	10162,
		40710	=>	10159,
		40711	=>	10157,
		40712	=>	10155,
		40713	=>	10153,
		40714	=>	10150,
		40715	=>	10148,
		40716	=>	10146,
		40717	=>	10143,
		40718	=>	10141,
		40719	=>	10139,
		40720	=>	10137,
		40721	=>	10134,
		40722	=>	10132,
		40723	=>	10130,
		40724	=>	10128,
		40725	=>	10125,
		40726	=>	10123,
		40727	=>	10121,
		40728	=>	10118,
		40729	=>	10116,
		40730	=>	10114,
		40731	=>	10112,
		40732	=>	10109,
		40733	=>	10107,
		40734	=>	10105,
		40735	=>	10103,
		40736	=>	10100,
		40737	=>	10098,
		40738	=>	10096,
		40739	=>	10093,
		40740	=>	10091,
		40741	=>	10089,
		40742	=>	10087,
		40743	=>	10084,
		40744	=>	10082,
		40745	=>	10080,
		40746	=>	10078,
		40747	=>	10075,
		40748	=>	10073,
		40749	=>	10071,
		40750	=>	10069,
		40751	=>	10066,
		40752	=>	10064,
		40753	=>	10062,
		40754	=>	10059,
		40755	=>	10057,
		40756	=>	10055,
		40757	=>	10053,
		40758	=>	10050,
		40759	=>	10048,
		40760	=>	10046,
		40761	=>	10044,
		40762	=>	10041,
		40763	=>	10039,
		40764	=>	10037,
		40765	=>	10035,
		40766	=>	10032,
		40767	=>	10030,
		40768	=>	10028,
		40769	=>	10026,
		40770	=>	10023,
		40771	=>	10021,
		40772	=>	10019,
		40773	=>	10016,
		40774	=>	10014,
		40775	=>	10012,
		40776	=>	10010,
		40777	=>	10007,
		40778	=>	10005,
		40779	=>	10003,
		40780	=>	10001,
		40781	=>	9998,
		40782	=>	9996,
		40783	=>	9994,
		40784	=>	9992,
		40785	=>	9989,
		40786	=>	9987,
		40787	=>	9985,
		40788	=>	9983,
		40789	=>	9980,
		40790	=>	9978,
		40791	=>	9976,
		40792	=>	9974,
		40793	=>	9971,
		40794	=>	9969,
		40795	=>	9967,
		40796	=>	9965,
		40797	=>	9962,
		40798	=>	9960,
		40799	=>	9958,
		40800	=>	9956,
		40801	=>	9953,
		40802	=>	9951,
		40803	=>	9949,
		40804	=>	9946,
		40805	=>	9944,
		40806	=>	9942,
		40807	=>	9940,
		40808	=>	9937,
		40809	=>	9935,
		40810	=>	9933,
		40811	=>	9931,
		40812	=>	9928,
		40813	=>	9926,
		40814	=>	9924,
		40815	=>	9922,
		40816	=>	9919,
		40817	=>	9917,
		40818	=>	9915,
		40819	=>	9913,
		40820	=>	9910,
		40821	=>	9908,
		40822	=>	9906,
		40823	=>	9904,
		40824	=>	9901,
		40825	=>	9899,
		40826	=>	9897,
		40827	=>	9895,
		40828	=>	9892,
		40829	=>	9890,
		40830	=>	9888,
		40831	=>	9886,
		40832	=>	9883,
		40833	=>	9881,
		40834	=>	9879,
		40835	=>	9877,
		40836	=>	9874,
		40837	=>	9872,
		40838	=>	9870,
		40839	=>	9868,
		40840	=>	9865,
		40841	=>	9863,
		40842	=>	9861,
		40843	=>	9859,
		40844	=>	9856,
		40845	=>	9854,
		40846	=>	9852,
		40847	=>	9850,
		40848	=>	9848,
		40849	=>	9845,
		40850	=>	9843,
		40851	=>	9841,
		40852	=>	9839,
		40853	=>	9836,
		40854	=>	9834,
		40855	=>	9832,
		40856	=>	9830,
		40857	=>	9827,
		40858	=>	9825,
		40859	=>	9823,
		40860	=>	9821,
		40861	=>	9818,
		40862	=>	9816,
		40863	=>	9814,
		40864	=>	9812,
		40865	=>	9809,
		40866	=>	9807,
		40867	=>	9805,
		40868	=>	9803,
		40869	=>	9800,
		40870	=>	9798,
		40871	=>	9796,
		40872	=>	9794,
		40873	=>	9791,
		40874	=>	9789,
		40875	=>	9787,
		40876	=>	9785,
		40877	=>	9782,
		40878	=>	9780,
		40879	=>	9778,
		40880	=>	9776,
		40881	=>	9774,
		40882	=>	9771,
		40883	=>	9769,
		40884	=>	9767,
		40885	=>	9765,
		40886	=>	9762,
		40887	=>	9760,
		40888	=>	9758,
		40889	=>	9756,
		40890	=>	9753,
		40891	=>	9751,
		40892	=>	9749,
		40893	=>	9747,
		40894	=>	9744,
		40895	=>	9742,
		40896	=>	9740,
		40897	=>	9738,
		40898	=>	9736,
		40899	=>	9733,
		40900	=>	9731,
		40901	=>	9729,
		40902	=>	9727,
		40903	=>	9724,
		40904	=>	9722,
		40905	=>	9720,
		40906	=>	9718,
		40907	=>	9715,
		40908	=>	9713,
		40909	=>	9711,
		40910	=>	9709,
		40911	=>	9706,
		40912	=>	9704,
		40913	=>	9702,
		40914	=>	9700,
		40915	=>	9698,
		40916	=>	9695,
		40917	=>	9693,
		40918	=>	9691,
		40919	=>	9689,
		40920	=>	9686,
		40921	=>	9684,
		40922	=>	9682,
		40923	=>	9680,
		40924	=>	9677,
		40925	=>	9675,
		40926	=>	9673,
		40927	=>	9671,
		40928	=>	9669,
		40929	=>	9666,
		40930	=>	9664,
		40931	=>	9662,
		40932	=>	9660,
		40933	=>	9657,
		40934	=>	9655,
		40935	=>	9653,
		40936	=>	9651,
		40937	=>	9649,
		40938	=>	9646,
		40939	=>	9644,
		40940	=>	9642,
		40941	=>	9640,
		40942	=>	9637,
		40943	=>	9635,
		40944	=>	9633,
		40945	=>	9631,
		40946	=>	9628,
		40947	=>	9626,
		40948	=>	9624,
		40949	=>	9622,
		40950	=>	9620,
		40951	=>	9617,
		40952	=>	9615,
		40953	=>	9613,
		40954	=>	9611,
		40955	=>	9608,
		40956	=>	9606,
		40957	=>	9604,
		40958	=>	9602,
		40959	=>	9600,
		40960	=>	9597,
		40961	=>	9595,
		40962	=>	9593,
		40963	=>	9591,
		40964	=>	9588,
		40965	=>	9586,
		40966	=>	9584,
		40967	=>	9582,
		40968	=>	9580,
		40969	=>	9577,
		40970	=>	9575,
		40971	=>	9573,
		40972	=>	9571,
		40973	=>	9569,
		40974	=>	9566,
		40975	=>	9564,
		40976	=>	9562,
		40977	=>	9560,
		40978	=>	9557,
		40979	=>	9555,
		40980	=>	9553,
		40981	=>	9551,
		40982	=>	9549,
		40983	=>	9546,
		40984	=>	9544,
		40985	=>	9542,
		40986	=>	9540,
		40987	=>	9537,
		40988	=>	9535,
		40989	=>	9533,
		40990	=>	9531,
		40991	=>	9529,
		40992	=>	9526,
		40993	=>	9524,
		40994	=>	9522,
		40995	=>	9520,
		40996	=>	9518,
		40997	=>	9515,
		40998	=>	9513,
		40999	=>	9511,
		41000	=>	9509,
		41001	=>	9506,
		41002	=>	9504,
		41003	=>	9502,
		41004	=>	9500,
		41005	=>	9498,
		41006	=>	9495,
		41007	=>	9493,
		41008	=>	9491,
		41009	=>	9489,
		41010	=>	9487,
		41011	=>	9484,
		41012	=>	9482,
		41013	=>	9480,
		41014	=>	9478,
		41015	=>	9476,
		41016	=>	9473,
		41017	=>	9471,
		41018	=>	9469,
		41019	=>	9467,
		41020	=>	9464,
		41021	=>	9462,
		41022	=>	9460,
		41023	=>	9458,
		41024	=>	9456,
		41025	=>	9453,
		41026	=>	9451,
		41027	=>	9449,
		41028	=>	9447,
		41029	=>	9445,
		41030	=>	9442,
		41031	=>	9440,
		41032	=>	9438,
		41033	=>	9436,
		41034	=>	9434,
		41035	=>	9431,
		41036	=>	9429,
		41037	=>	9427,
		41038	=>	9425,
		41039	=>	9423,
		41040	=>	9420,
		41041	=>	9418,
		41042	=>	9416,
		41043	=>	9414,
		41044	=>	9412,
		41045	=>	9409,
		41046	=>	9407,
		41047	=>	9405,
		41048	=>	9403,
		41049	=>	9401,
		41050	=>	9398,
		41051	=>	9396,
		41052	=>	9394,
		41053	=>	9392,
		41054	=>	9390,
		41055	=>	9387,
		41056	=>	9385,
		41057	=>	9383,
		41058	=>	9381,
		41059	=>	9379,
		41060	=>	9376,
		41061	=>	9374,
		41062	=>	9372,
		41063	=>	9370,
		41064	=>	9368,
		41065	=>	9365,
		41066	=>	9363,
		41067	=>	9361,
		41068	=>	9359,
		41069	=>	9357,
		41070	=>	9354,
		41071	=>	9352,
		41072	=>	9350,
		41073	=>	9348,
		41074	=>	9346,
		41075	=>	9343,
		41076	=>	9341,
		41077	=>	9339,
		41078	=>	9337,
		41079	=>	9335,
		41080	=>	9332,
		41081	=>	9330,
		41082	=>	9328,
		41083	=>	9326,
		41084	=>	9324,
		41085	=>	9321,
		41086	=>	9319,
		41087	=>	9317,
		41088	=>	9315,
		41089	=>	9313,
		41090	=>	9310,
		41091	=>	9308,
		41092	=>	9306,
		41093	=>	9304,
		41094	=>	9302,
		41095	=>	9299,
		41096	=>	9297,
		41097	=>	9295,
		41098	=>	9293,
		41099	=>	9291,
		41100	=>	9288,
		41101	=>	9286,
		41102	=>	9284,
		41103	=>	9282,
		41104	=>	9280,
		41105	=>	9278,
		41106	=>	9275,
		41107	=>	9273,
		41108	=>	9271,
		41109	=>	9269,
		41110	=>	9267,
		41111	=>	9264,
		41112	=>	9262,
		41113	=>	9260,
		41114	=>	9258,
		41115	=>	9256,
		41116	=>	9253,
		41117	=>	9251,
		41118	=>	9249,
		41119	=>	9247,
		41120	=>	9245,
		41121	=>	9243,
		41122	=>	9240,
		41123	=>	9238,
		41124	=>	9236,
		41125	=>	9234,
		41126	=>	9232,
		41127	=>	9229,
		41128	=>	9227,
		41129	=>	9225,
		41130	=>	9223,
		41131	=>	9221,
		41132	=>	9218,
		41133	=>	9216,
		41134	=>	9214,
		41135	=>	9212,
		41136	=>	9210,
		41137	=>	9208,
		41138	=>	9205,
		41139	=>	9203,
		41140	=>	9201,
		41141	=>	9199,
		41142	=>	9197,
		41143	=>	9194,
		41144	=>	9192,
		41145	=>	9190,
		41146	=>	9188,
		41147	=>	9186,
		41148	=>	9184,
		41149	=>	9181,
		41150	=>	9179,
		41151	=>	9177,
		41152	=>	9175,
		41153	=>	9173,
		41154	=>	9170,
		41155	=>	9168,
		41156	=>	9166,
		41157	=>	9164,
		41158	=>	9162,
		41159	=>	9160,
		41160	=>	9157,
		41161	=>	9155,
		41162	=>	9153,
		41163	=>	9151,
		41164	=>	9149,
		41165	=>	9146,
		41166	=>	9144,
		41167	=>	9142,
		41168	=>	9140,
		41169	=>	9138,
		41170	=>	9136,
		41171	=>	9133,
		41172	=>	9131,
		41173	=>	9129,
		41174	=>	9127,
		41175	=>	9125,
		41176	=>	9123,
		41177	=>	9120,
		41178	=>	9118,
		41179	=>	9116,
		41180	=>	9114,
		41181	=>	9112,
		41182	=>	9110,
		41183	=>	9107,
		41184	=>	9105,
		41185	=>	9103,
		41186	=>	9101,
		41187	=>	9099,
		41188	=>	9096,
		41189	=>	9094,
		41190	=>	9092,
		41191	=>	9090,
		41192	=>	9088,
		41193	=>	9086,
		41194	=>	9083,
		41195	=>	9081,
		41196	=>	9079,
		41197	=>	9077,
		41198	=>	9075,
		41199	=>	9073,
		41200	=>	9070,
		41201	=>	9068,
		41202	=>	9066,
		41203	=>	9064,
		41204	=>	9062,
		41205	=>	9060,
		41206	=>	9057,
		41207	=>	9055,
		41208	=>	9053,
		41209	=>	9051,
		41210	=>	9049,
		41211	=>	9047,
		41212	=>	9044,
		41213	=>	9042,
		41214	=>	9040,
		41215	=>	9038,
		41216	=>	9036,
		41217	=>	9034,
		41218	=>	9031,
		41219	=>	9029,
		41220	=>	9027,
		41221	=>	9025,
		41222	=>	9023,
		41223	=>	9021,
		41224	=>	9018,
		41225	=>	9016,
		41226	=>	9014,
		41227	=>	9012,
		41228	=>	9010,
		41229	=>	9008,
		41230	=>	9005,
		41231	=>	9003,
		41232	=>	9001,
		41233	=>	8999,
		41234	=>	8997,
		41235	=>	8995,
		41236	=>	8992,
		41237	=>	8990,
		41238	=>	8988,
		41239	=>	8986,
		41240	=>	8984,
		41241	=>	8982,
		41242	=>	8979,
		41243	=>	8977,
		41244	=>	8975,
		41245	=>	8973,
		41246	=>	8971,
		41247	=>	8969,
		41248	=>	8967,
		41249	=>	8964,
		41250	=>	8962,
		41251	=>	8960,
		41252	=>	8958,
		41253	=>	8956,
		41254	=>	8954,
		41255	=>	8951,
		41256	=>	8949,
		41257	=>	8947,
		41258	=>	8945,
		41259	=>	8943,
		41260	=>	8941,
		41261	=>	8938,
		41262	=>	8936,
		41263	=>	8934,
		41264	=>	8932,
		41265	=>	8930,
		41266	=>	8928,
		41267	=>	8926,
		41268	=>	8923,
		41269	=>	8921,
		41270	=>	8919,
		41271	=>	8917,
		41272	=>	8915,
		41273	=>	8913,
		41274	=>	8910,
		41275	=>	8908,
		41276	=>	8906,
		41277	=>	8904,
		41278	=>	8902,
		41279	=>	8900,
		41280	=>	8898,
		41281	=>	8895,
		41282	=>	8893,
		41283	=>	8891,
		41284	=>	8889,
		41285	=>	8887,
		41286	=>	8885,
		41287	=>	8882,
		41288	=>	8880,
		41289	=>	8878,
		41290	=>	8876,
		41291	=>	8874,
		41292	=>	8872,
		41293	=>	8870,
		41294	=>	8867,
		41295	=>	8865,
		41296	=>	8863,
		41297	=>	8861,
		41298	=>	8859,
		41299	=>	8857,
		41300	=>	8855,
		41301	=>	8852,
		41302	=>	8850,
		41303	=>	8848,
		41304	=>	8846,
		41305	=>	8844,
		41306	=>	8842,
		41307	=>	8840,
		41308	=>	8837,
		41309	=>	8835,
		41310	=>	8833,
		41311	=>	8831,
		41312	=>	8829,
		41313	=>	8827,
		41314	=>	8824,
		41315	=>	8822,
		41316	=>	8820,
		41317	=>	8818,
		41318	=>	8816,
		41319	=>	8814,
		41320	=>	8812,
		41321	=>	8809,
		41322	=>	8807,
		41323	=>	8805,
		41324	=>	8803,
		41325	=>	8801,
		41326	=>	8799,
		41327	=>	8797,
		41328	=>	8794,
		41329	=>	8792,
		41330	=>	8790,
		41331	=>	8788,
		41332	=>	8786,
		41333	=>	8784,
		41334	=>	8782,
		41335	=>	8780,
		41336	=>	8777,
		41337	=>	8775,
		41338	=>	8773,
		41339	=>	8771,
		41340	=>	8769,
		41341	=>	8767,
		41342	=>	8765,
		41343	=>	8762,
		41344	=>	8760,
		41345	=>	8758,
		41346	=>	8756,
		41347	=>	8754,
		41348	=>	8752,
		41349	=>	8750,
		41350	=>	8747,
		41351	=>	8745,
		41352	=>	8743,
		41353	=>	8741,
		41354	=>	8739,
		41355	=>	8737,
		41356	=>	8735,
		41357	=>	8732,
		41358	=>	8730,
		41359	=>	8728,
		41360	=>	8726,
		41361	=>	8724,
		41362	=>	8722,
		41363	=>	8720,
		41364	=>	8718,
		41365	=>	8715,
		41366	=>	8713,
		41367	=>	8711,
		41368	=>	8709,
		41369	=>	8707,
		41370	=>	8705,
		41371	=>	8703,
		41372	=>	8700,
		41373	=>	8698,
		41374	=>	8696,
		41375	=>	8694,
		41376	=>	8692,
		41377	=>	8690,
		41378	=>	8688,
		41379	=>	8686,
		41380	=>	8683,
		41381	=>	8681,
		41382	=>	8679,
		41383	=>	8677,
		41384	=>	8675,
		41385	=>	8673,
		41386	=>	8671,
		41387	=>	8669,
		41388	=>	8666,
		41389	=>	8664,
		41390	=>	8662,
		41391	=>	8660,
		41392	=>	8658,
		41393	=>	8656,
		41394	=>	8654,
		41395	=>	8651,
		41396	=>	8649,
		41397	=>	8647,
		41398	=>	8645,
		41399	=>	8643,
		41400	=>	8641,
		41401	=>	8639,
		41402	=>	8637,
		41403	=>	8634,
		41404	=>	8632,
		41405	=>	8630,
		41406	=>	8628,
		41407	=>	8626,
		41408	=>	8624,
		41409	=>	8622,
		41410	=>	8620,
		41411	=>	8617,
		41412	=>	8615,
		41413	=>	8613,
		41414	=>	8611,
		41415	=>	8609,
		41416	=>	8607,
		41417	=>	8605,
		41418	=>	8603,
		41419	=>	8601,
		41420	=>	8598,
		41421	=>	8596,
		41422	=>	8594,
		41423	=>	8592,
		41424	=>	8590,
		41425	=>	8588,
		41426	=>	8586,
		41427	=>	8584,
		41428	=>	8581,
		41429	=>	8579,
		41430	=>	8577,
		41431	=>	8575,
		41432	=>	8573,
		41433	=>	8571,
		41434	=>	8569,
		41435	=>	8567,
		41436	=>	8564,
		41437	=>	8562,
		41438	=>	8560,
		41439	=>	8558,
		41440	=>	8556,
		41441	=>	8554,
		41442	=>	8552,
		41443	=>	8550,
		41444	=>	8548,
		41445	=>	8545,
		41446	=>	8543,
		41447	=>	8541,
		41448	=>	8539,
		41449	=>	8537,
		41450	=>	8535,
		41451	=>	8533,
		41452	=>	8531,
		41453	=>	8529,
		41454	=>	8526,
		41455	=>	8524,
		41456	=>	8522,
		41457	=>	8520,
		41458	=>	8518,
		41459	=>	8516,
		41460	=>	8514,
		41461	=>	8512,
		41462	=>	8509,
		41463	=>	8507,
		41464	=>	8505,
		41465	=>	8503,
		41466	=>	8501,
		41467	=>	8499,
		41468	=>	8497,
		41469	=>	8495,
		41470	=>	8493,
		41471	=>	8490,
		41472	=>	8488,
		41473	=>	8486,
		41474	=>	8484,
		41475	=>	8482,
		41476	=>	8480,
		41477	=>	8478,
		41478	=>	8476,
		41479	=>	8474,
		41480	=>	8472,
		41481	=>	8469,
		41482	=>	8467,
		41483	=>	8465,
		41484	=>	8463,
		41485	=>	8461,
		41486	=>	8459,
		41487	=>	8457,
		41488	=>	8455,
		41489	=>	8453,
		41490	=>	8450,
		41491	=>	8448,
		41492	=>	8446,
		41493	=>	8444,
		41494	=>	8442,
		41495	=>	8440,
		41496	=>	8438,
		41497	=>	8436,
		41498	=>	8434,
		41499	=>	8432,
		41500	=>	8429,
		41501	=>	8427,
		41502	=>	8425,
		41503	=>	8423,
		41504	=>	8421,
		41505	=>	8419,
		41506	=>	8417,
		41507	=>	8415,
		41508	=>	8413,
		41509	=>	8410,
		41510	=>	8408,
		41511	=>	8406,
		41512	=>	8404,
		41513	=>	8402,
		41514	=>	8400,
		41515	=>	8398,
		41516	=>	8396,
		41517	=>	8394,
		41518	=>	8392,
		41519	=>	8389,
		41520	=>	8387,
		41521	=>	8385,
		41522	=>	8383,
		41523	=>	8381,
		41524	=>	8379,
		41525	=>	8377,
		41526	=>	8375,
		41527	=>	8373,
		41528	=>	8371,
		41529	=>	8368,
		41530	=>	8366,
		41531	=>	8364,
		41532	=>	8362,
		41533	=>	8360,
		41534	=>	8358,
		41535	=>	8356,
		41536	=>	8354,
		41537	=>	8352,
		41538	=>	8350,
		41539	=>	8348,
		41540	=>	8345,
		41541	=>	8343,
		41542	=>	8341,
		41543	=>	8339,
		41544	=>	8337,
		41545	=>	8335,
		41546	=>	8333,
		41547	=>	8331,
		41548	=>	8329,
		41549	=>	8327,
		41550	=>	8325,
		41551	=>	8322,
		41552	=>	8320,
		41553	=>	8318,
		41554	=>	8316,
		41555	=>	8314,
		41556	=>	8312,
		41557	=>	8310,
		41558	=>	8308,
		41559	=>	8306,
		41560	=>	8304,
		41561	=>	8302,
		41562	=>	8299,
		41563	=>	8297,
		41564	=>	8295,
		41565	=>	8293,
		41566	=>	8291,
		41567	=>	8289,
		41568	=>	8287,
		41569	=>	8285,
		41570	=>	8283,
		41571	=>	8281,
		41572	=>	8279,
		41573	=>	8276,
		41574	=>	8274,
		41575	=>	8272,
		41576	=>	8270,
		41577	=>	8268,
		41578	=>	8266,
		41579	=>	8264,
		41580	=>	8262,
		41581	=>	8260,
		41582	=>	8258,
		41583	=>	8256,
		41584	=>	8253,
		41585	=>	8251,
		41586	=>	8249,
		41587	=>	8247,
		41588	=>	8245,
		41589	=>	8243,
		41590	=>	8241,
		41591	=>	8239,
		41592	=>	8237,
		41593	=>	8235,
		41594	=>	8233,
		41595	=>	8231,
		41596	=>	8228,
		41597	=>	8226,
		41598	=>	8224,
		41599	=>	8222,
		41600	=>	8220,
		41601	=>	8218,
		41602	=>	8216,
		41603	=>	8214,
		41604	=>	8212,
		41605	=>	8210,
		41606	=>	8208,
		41607	=>	8206,
		41608	=>	8204,
		41609	=>	8201,
		41610	=>	8199,
		41611	=>	8197,
		41612	=>	8195,
		41613	=>	8193,
		41614	=>	8191,
		41615	=>	8189,
		41616	=>	8187,
		41617	=>	8185,
		41618	=>	8183,
		41619	=>	8181,
		41620	=>	8179,
		41621	=>	8177,
		41622	=>	8174,
		41623	=>	8172,
		41624	=>	8170,
		41625	=>	8168,
		41626	=>	8166,
		41627	=>	8164,
		41628	=>	8162,
		41629	=>	8160,
		41630	=>	8158,
		41631	=>	8156,
		41632	=>	8154,
		41633	=>	8152,
		41634	=>	8150,
		41635	=>	8147,
		41636	=>	8145,
		41637	=>	8143,
		41638	=>	8141,
		41639	=>	8139,
		41640	=>	8137,
		41641	=>	8135,
		41642	=>	8133,
		41643	=>	8131,
		41644	=>	8129,
		41645	=>	8127,
		41646	=>	8125,
		41647	=>	8123,
		41648	=>	8121,
		41649	=>	8118,
		41650	=>	8116,
		41651	=>	8114,
		41652	=>	8112,
		41653	=>	8110,
		41654	=>	8108,
		41655	=>	8106,
		41656	=>	8104,
		41657	=>	8102,
		41658	=>	8100,
		41659	=>	8098,
		41660	=>	8096,
		41661	=>	8094,
		41662	=>	8092,
		41663	=>	8090,
		41664	=>	8087,
		41665	=>	8085,
		41666	=>	8083,
		41667	=>	8081,
		41668	=>	8079,
		41669	=>	8077,
		41670	=>	8075,
		41671	=>	8073,
		41672	=>	8071,
		41673	=>	8069,
		41674	=>	8067,
		41675	=>	8065,
		41676	=>	8063,
		41677	=>	8061,
		41678	=>	8059,
		41679	=>	8056,
		41680	=>	8054,
		41681	=>	8052,
		41682	=>	8050,
		41683	=>	8048,
		41684	=>	8046,
		41685	=>	8044,
		41686	=>	8042,
		41687	=>	8040,
		41688	=>	8038,
		41689	=>	8036,
		41690	=>	8034,
		41691	=>	8032,
		41692	=>	8030,
		41693	=>	8028,
		41694	=>	8026,
		41695	=>	8023,
		41696	=>	8021,
		41697	=>	8019,
		41698	=>	8017,
		41699	=>	8015,
		41700	=>	8013,
		41701	=>	8011,
		41702	=>	8009,
		41703	=>	8007,
		41704	=>	8005,
		41705	=>	8003,
		41706	=>	8001,
		41707	=>	7999,
		41708	=>	7997,
		41709	=>	7995,
		41710	=>	7993,
		41711	=>	7991,
		41712	=>	7989,
		41713	=>	7986,
		41714	=>	7984,
		41715	=>	7982,
		41716	=>	7980,
		41717	=>	7978,
		41718	=>	7976,
		41719	=>	7974,
		41720	=>	7972,
		41721	=>	7970,
		41722	=>	7968,
		41723	=>	7966,
		41724	=>	7964,
		41725	=>	7962,
		41726	=>	7960,
		41727	=>	7958,
		41728	=>	7956,
		41729	=>	7954,
		41730	=>	7952,
		41731	=>	7950,
		41732	=>	7947,
		41733	=>	7945,
		41734	=>	7943,
		41735	=>	7941,
		41736	=>	7939,
		41737	=>	7937,
		41738	=>	7935,
		41739	=>	7933,
		41740	=>	7931,
		41741	=>	7929,
		41742	=>	7927,
		41743	=>	7925,
		41744	=>	7923,
		41745	=>	7921,
		41746	=>	7919,
		41747	=>	7917,
		41748	=>	7915,
		41749	=>	7913,
		41750	=>	7911,
		41751	=>	7909,
		41752	=>	7906,
		41753	=>	7904,
		41754	=>	7902,
		41755	=>	7900,
		41756	=>	7898,
		41757	=>	7896,
		41758	=>	7894,
		41759	=>	7892,
		41760	=>	7890,
		41761	=>	7888,
		41762	=>	7886,
		41763	=>	7884,
		41764	=>	7882,
		41765	=>	7880,
		41766	=>	7878,
		41767	=>	7876,
		41768	=>	7874,
		41769	=>	7872,
		41770	=>	7870,
		41771	=>	7868,
		41772	=>	7866,
		41773	=>	7864,
		41774	=>	7862,
		41775	=>	7859,
		41776	=>	7857,
		41777	=>	7855,
		41778	=>	7853,
		41779	=>	7851,
		41780	=>	7849,
		41781	=>	7847,
		41782	=>	7845,
		41783	=>	7843,
		41784	=>	7841,
		41785	=>	7839,
		41786	=>	7837,
		41787	=>	7835,
		41788	=>	7833,
		41789	=>	7831,
		41790	=>	7829,
		41791	=>	7827,
		41792	=>	7825,
		41793	=>	7823,
		41794	=>	7821,
		41795	=>	7819,
		41796	=>	7817,
		41797	=>	7815,
		41798	=>	7813,
		41799	=>	7811,
		41800	=>	7809,
		41801	=>	7806,
		41802	=>	7804,
		41803	=>	7802,
		41804	=>	7800,
		41805	=>	7798,
		41806	=>	7796,
		41807	=>	7794,
		41808	=>	7792,
		41809	=>	7790,
		41810	=>	7788,
		41811	=>	7786,
		41812	=>	7784,
		41813	=>	7782,
		41814	=>	7780,
		41815	=>	7778,
		41816	=>	7776,
		41817	=>	7774,
		41818	=>	7772,
		41819	=>	7770,
		41820	=>	7768,
		41821	=>	7766,
		41822	=>	7764,
		41823	=>	7762,
		41824	=>	7760,
		41825	=>	7758,
		41826	=>	7756,
		41827	=>	7754,
		41828	=>	7752,
		41829	=>	7750,
		41830	=>	7748,
		41831	=>	7746,
		41832	=>	7743,
		41833	=>	7741,
		41834	=>	7739,
		41835	=>	7737,
		41836	=>	7735,
		41837	=>	7733,
		41838	=>	7731,
		41839	=>	7729,
		41840	=>	7727,
		41841	=>	7725,
		41842	=>	7723,
		41843	=>	7721,
		41844	=>	7719,
		41845	=>	7717,
		41846	=>	7715,
		41847	=>	7713,
		41848	=>	7711,
		41849	=>	7709,
		41850	=>	7707,
		41851	=>	7705,
		41852	=>	7703,
		41853	=>	7701,
		41854	=>	7699,
		41855	=>	7697,
		41856	=>	7695,
		41857	=>	7693,
		41858	=>	7691,
		41859	=>	7689,
		41860	=>	7687,
		41861	=>	7685,
		41862	=>	7683,
		41863	=>	7681,
		41864	=>	7679,
		41865	=>	7677,
		41866	=>	7675,
		41867	=>	7673,
		41868	=>	7671,
		41869	=>	7669,
		41870	=>	7667,
		41871	=>	7665,
		41872	=>	7663,
		41873	=>	7661,
		41874	=>	7659,
		41875	=>	7656,
		41876	=>	7654,
		41877	=>	7652,
		41878	=>	7650,
		41879	=>	7648,
		41880	=>	7646,
		41881	=>	7644,
		41882	=>	7642,
		41883	=>	7640,
		41884	=>	7638,
		41885	=>	7636,
		41886	=>	7634,
		41887	=>	7632,
		41888	=>	7630,
		41889	=>	7628,
		41890	=>	7626,
		41891	=>	7624,
		41892	=>	7622,
		41893	=>	7620,
		41894	=>	7618,
		41895	=>	7616,
		41896	=>	7614,
		41897	=>	7612,
		41898	=>	7610,
		41899	=>	7608,
		41900	=>	7606,
		41901	=>	7604,
		41902	=>	7602,
		41903	=>	7600,
		41904	=>	7598,
		41905	=>	7596,
		41906	=>	7594,
		41907	=>	7592,
		41908	=>	7590,
		41909	=>	7588,
		41910	=>	7586,
		41911	=>	7584,
		41912	=>	7582,
		41913	=>	7580,
		41914	=>	7578,
		41915	=>	7576,
		41916	=>	7574,
		41917	=>	7572,
		41918	=>	7570,
		41919	=>	7568,
		41920	=>	7566,
		41921	=>	7564,
		41922	=>	7562,
		41923	=>	7560,
		41924	=>	7558,
		41925	=>	7556,
		41926	=>	7554,
		41927	=>	7552,
		41928	=>	7550,
		41929	=>	7548,
		41930	=>	7546,
		41931	=>	7544,
		41932	=>	7542,
		41933	=>	7540,
		41934	=>	7538,
		41935	=>	7536,
		41936	=>	7534,
		41937	=>	7532,
		41938	=>	7530,
		41939	=>	7528,
		41940	=>	7526,
		41941	=>	7524,
		41942	=>	7522,
		41943	=>	7520,
		41944	=>	7518,
		41945	=>	7516,
		41946	=>	7514,
		41947	=>	7512,
		41948	=>	7510,
		41949	=>	7508,
		41950	=>	7506,
		41951	=>	7504,
		41952	=>	7502,
		41953	=>	7500,
		41954	=>	7498,
		41955	=>	7496,
		41956	=>	7494,
		41957	=>	7492,
		41958	=>	7490,
		41959	=>	7488,
		41960	=>	7486,
		41961	=>	7484,
		41962	=>	7482,
		41963	=>	7480,
		41964	=>	7478,
		41965	=>	7476,
		41966	=>	7474,
		41967	=>	7472,
		41968	=>	7470,
		41969	=>	7468,
		41970	=>	7466,
		41971	=>	7464,
		41972	=>	7462,
		41973	=>	7460,
		41974	=>	7458,
		41975	=>	7456,
		41976	=>	7454,
		41977	=>	7452,
		41978	=>	7450,
		41979	=>	7448,
		41980	=>	7446,
		41981	=>	7444,
		41982	=>	7442,
		41983	=>	7440,
		41984	=>	7438,
		41985	=>	7436,
		41986	=>	7434,
		41987	=>	7432,
		41988	=>	7430,
		41989	=>	7428,
		41990	=>	7426,
		41991	=>	7424,
		41992	=>	7422,
		41993	=>	7420,
		41994	=>	7418,
		41995	=>	7416,
		41996	=>	7414,
		41997	=>	7412,
		41998	=>	7410,
		41999	=>	7408,
		42000	=>	7406,
		42001	=>	7404,
		42002	=>	7402,
		42003	=>	7400,
		42004	=>	7398,
		42005	=>	7396,
		42006	=>	7394,
		42007	=>	7392,
		42008	=>	7390,
		42009	=>	7388,
		42010	=>	7386,
		42011	=>	7384,
		42012	=>	7382,
		42013	=>	7380,
		42014	=>	7378,
		42015	=>	7376,
		42016	=>	7374,
		42017	=>	7372,
		42018	=>	7370,
		42019	=>	7368,
		42020	=>	7366,
		42021	=>	7364,
		42022	=>	7362,
		42023	=>	7360,
		42024	=>	7358,
		42025	=>	7356,
		42026	=>	7354,
		42027	=>	7352,
		42028	=>	7350,
		42029	=>	7348,
		42030	=>	7346,
		42031	=>	7344,
		42032	=>	7342,
		42033	=>	7341,
		42034	=>	7339,
		42035	=>	7337,
		42036	=>	7335,
		42037	=>	7333,
		42038	=>	7331,
		42039	=>	7329,
		42040	=>	7327,
		42041	=>	7325,
		42042	=>	7323,
		42043	=>	7321,
		42044	=>	7319,
		42045	=>	7317,
		42046	=>	7315,
		42047	=>	7313,
		42048	=>	7311,
		42049	=>	7309,
		42050	=>	7307,
		42051	=>	7305,
		42052	=>	7303,
		42053	=>	7301,
		42054	=>	7299,
		42055	=>	7297,
		42056	=>	7295,
		42057	=>	7293,
		42058	=>	7291,
		42059	=>	7289,
		42060	=>	7287,
		42061	=>	7285,
		42062	=>	7283,
		42063	=>	7281,
		42064	=>	7279,
		42065	=>	7277,
		42066	=>	7275,
		42067	=>	7273,
		42068	=>	7271,
		42069	=>	7269,
		42070	=>	7267,
		42071	=>	7265,
		42072	=>	7263,
		42073	=>	7261,
		42074	=>	7259,
		42075	=>	7257,
		42076	=>	7256,
		42077	=>	7254,
		42078	=>	7252,
		42079	=>	7250,
		42080	=>	7248,
		42081	=>	7246,
		42082	=>	7244,
		42083	=>	7242,
		42084	=>	7240,
		42085	=>	7238,
		42086	=>	7236,
		42087	=>	7234,
		42088	=>	7232,
		42089	=>	7230,
		42090	=>	7228,
		42091	=>	7226,
		42092	=>	7224,
		42093	=>	7222,
		42094	=>	7220,
		42095	=>	7218,
		42096	=>	7216,
		42097	=>	7214,
		42098	=>	7212,
		42099	=>	7210,
		42100	=>	7208,
		42101	=>	7206,
		42102	=>	7204,
		42103	=>	7202,
		42104	=>	7200,
		42105	=>	7198,
		42106	=>	7196,
		42107	=>	7195,
		42108	=>	7193,
		42109	=>	7191,
		42110	=>	7189,
		42111	=>	7187,
		42112	=>	7185,
		42113	=>	7183,
		42114	=>	7181,
		42115	=>	7179,
		42116	=>	7177,
		42117	=>	7175,
		42118	=>	7173,
		42119	=>	7171,
		42120	=>	7169,
		42121	=>	7167,
		42122	=>	7165,
		42123	=>	7163,
		42124	=>	7161,
		42125	=>	7159,
		42126	=>	7157,
		42127	=>	7155,
		42128	=>	7153,
		42129	=>	7151,
		42130	=>	7149,
		42131	=>	7147,
		42132	=>	7145,
		42133	=>	7144,
		42134	=>	7142,
		42135	=>	7140,
		42136	=>	7138,
		42137	=>	7136,
		42138	=>	7134,
		42139	=>	7132,
		42140	=>	7130,
		42141	=>	7128,
		42142	=>	7126,
		42143	=>	7124,
		42144	=>	7122,
		42145	=>	7120,
		42146	=>	7118,
		42147	=>	7116,
		42148	=>	7114,
		42149	=>	7112,
		42150	=>	7110,
		42151	=>	7108,
		42152	=>	7106,
		42153	=>	7104,
		42154	=>	7102,
		42155	=>	7101,
		42156	=>	7099,
		42157	=>	7097,
		42158	=>	7095,
		42159	=>	7093,
		42160	=>	7091,
		42161	=>	7089,
		42162	=>	7087,
		42163	=>	7085,
		42164	=>	7083,
		42165	=>	7081,
		42166	=>	7079,
		42167	=>	7077,
		42168	=>	7075,
		42169	=>	7073,
		42170	=>	7071,
		42171	=>	7069,
		42172	=>	7067,
		42173	=>	7065,
		42174	=>	7063,
		42175	=>	7061,
		42176	=>	7060,
		42177	=>	7058,
		42178	=>	7056,
		42179	=>	7054,
		42180	=>	7052,
		42181	=>	7050,
		42182	=>	7048,
		42183	=>	7046,
		42184	=>	7044,
		42185	=>	7042,
		42186	=>	7040,
		42187	=>	7038,
		42188	=>	7036,
		42189	=>	7034,
		42190	=>	7032,
		42191	=>	7030,
		42192	=>	7028,
		42193	=>	7026,
		42194	=>	7025,
		42195	=>	7023,
		42196	=>	7021,
		42197	=>	7019,
		42198	=>	7017,
		42199	=>	7015,
		42200	=>	7013,
		42201	=>	7011,
		42202	=>	7009,
		42203	=>	7007,
		42204	=>	7005,
		42205	=>	7003,
		42206	=>	7001,
		42207	=>	6999,
		42208	=>	6997,
		42209	=>	6995,
		42210	=>	6993,
		42211	=>	6992,
		42212	=>	6990,
		42213	=>	6988,
		42214	=>	6986,
		42215	=>	6984,
		42216	=>	6982,
		42217	=>	6980,
		42218	=>	6978,
		42219	=>	6976,
		42220	=>	6974,
		42221	=>	6972,
		42222	=>	6970,
		42223	=>	6968,
		42224	=>	6966,
		42225	=>	6964,
		42226	=>	6962,
		42227	=>	6961,
		42228	=>	6959,
		42229	=>	6957,
		42230	=>	6955,
		42231	=>	6953,
		42232	=>	6951,
		42233	=>	6949,
		42234	=>	6947,
		42235	=>	6945,
		42236	=>	6943,
		42237	=>	6941,
		42238	=>	6939,
		42239	=>	6937,
		42240	=>	6935,
		42241	=>	6933,
		42242	=>	6931,
		42243	=>	6930,
		42244	=>	6928,
		42245	=>	6926,
		42246	=>	6924,
		42247	=>	6922,
		42248	=>	6920,
		42249	=>	6918,
		42250	=>	6916,
		42251	=>	6914,
		42252	=>	6912,
		42253	=>	6910,
		42254	=>	6908,
		42255	=>	6906,
		42256	=>	6904,
		42257	=>	6903,
		42258	=>	6901,
		42259	=>	6899,
		42260	=>	6897,
		42261	=>	6895,
		42262	=>	6893,
		42263	=>	6891,
		42264	=>	6889,
		42265	=>	6887,
		42266	=>	6885,
		42267	=>	6883,
		42268	=>	6881,
		42269	=>	6879,
		42270	=>	6877,
		42271	=>	6876,
		42272	=>	6874,
		42273	=>	6872,
		42274	=>	6870,
		42275	=>	6868,
		42276	=>	6866,
		42277	=>	6864,
		42278	=>	6862,
		42279	=>	6860,
		42280	=>	6858,
		42281	=>	6856,
		42282	=>	6854,
		42283	=>	6852,
		42284	=>	6851,
		42285	=>	6849,
		42286	=>	6847,
		42287	=>	6845,
		42288	=>	6843,
		42289	=>	6841,
		42290	=>	6839,
		42291	=>	6837,
		42292	=>	6835,
		42293	=>	6833,
		42294	=>	6831,
		42295	=>	6829,
		42296	=>	6827,
		42297	=>	6826,
		42298	=>	6824,
		42299	=>	6822,
		42300	=>	6820,
		42301	=>	6818,
		42302	=>	6816,
		42303	=>	6814,
		42304	=>	6812,
		42305	=>	6810,
		42306	=>	6808,
		42307	=>	6806,
		42308	=>	6804,
		42309	=>	6803,
		42310	=>	6801,
		42311	=>	6799,
		42312	=>	6797,
		42313	=>	6795,
		42314	=>	6793,
		42315	=>	6791,
		42316	=>	6789,
		42317	=>	6787,
		42318	=>	6785,
		42319	=>	6783,
		42320	=>	6781,
		42321	=>	6780,
		42322	=>	6778,
		42323	=>	6776,
		42324	=>	6774,
		42325	=>	6772,
		42326	=>	6770,
		42327	=>	6768,
		42328	=>	6766,
		42329	=>	6764,
		42330	=>	6762,
		42331	=>	6760,
		42332	=>	6759,
		42333	=>	6757,
		42334	=>	6755,
		42335	=>	6753,
		42336	=>	6751,
		42337	=>	6749,
		42338	=>	6747,
		42339	=>	6745,
		42340	=>	6743,
		42341	=>	6741,
		42342	=>	6739,
		42343	=>	6738,
		42344	=>	6736,
		42345	=>	6734,
		42346	=>	6732,
		42347	=>	6730,
		42348	=>	6728,
		42349	=>	6726,
		42350	=>	6724,
		42351	=>	6722,
		42352	=>	6720,
		42353	=>	6718,
		42354	=>	6717,
		42355	=>	6715,
		42356	=>	6713,
		42357	=>	6711,
		42358	=>	6709,
		42359	=>	6707,
		42360	=>	6705,
		42361	=>	6703,
		42362	=>	6701,
		42363	=>	6699,
		42364	=>	6698,
		42365	=>	6696,
		42366	=>	6694,
		42367	=>	6692,
		42368	=>	6690,
		42369	=>	6688,
		42370	=>	6686,
		42371	=>	6684,
		42372	=>	6682,
		42373	=>	6680,
		42374	=>	6679,
		42375	=>	6677,
		42376	=>	6675,
		42377	=>	6673,
		42378	=>	6671,
		42379	=>	6669,
		42380	=>	6667,
		42381	=>	6665,
		42382	=>	6663,
		42383	=>	6661,
		42384	=>	6660,
		42385	=>	6658,
		42386	=>	6656,
		42387	=>	6654,
		42388	=>	6652,
		42389	=>	6650,
		42390	=>	6648,
		42391	=>	6646,
		42392	=>	6644,
		42393	=>	6642,
		42394	=>	6641,
		42395	=>	6639,
		42396	=>	6637,
		42397	=>	6635,
		42398	=>	6633,
		42399	=>	6631,
		42400	=>	6629,
		42401	=>	6627,
		42402	=>	6625,
		42403	=>	6623,
		42404	=>	6622,
		42405	=>	6620,
		42406	=>	6618,
		42407	=>	6616,
		42408	=>	6614,
		42409	=>	6612,
		42410	=>	6610,
		42411	=>	6608,
		42412	=>	6606,
		42413	=>	6605,
		42414	=>	6603,
		42415	=>	6601,
		42416	=>	6599,
		42417	=>	6597,
		42418	=>	6595,
		42419	=>	6593,
		42420	=>	6591,
		42421	=>	6589,
		42422	=>	6588,
		42423	=>	6586,
		42424	=>	6584,
		42425	=>	6582,
		42426	=>	6580,
		42427	=>	6578,
		42428	=>	6576,
		42429	=>	6574,
		42430	=>	6572,
		42431	=>	6571,
		42432	=>	6569,
		42433	=>	6567,
		42434	=>	6565,
		42435	=>	6563,
		42436	=>	6561,
		42437	=>	6559,
		42438	=>	6557,
		42439	=>	6555,
		42440	=>	6554,
		42441	=>	6552,
		42442	=>	6550,
		42443	=>	6548,
		42444	=>	6546,
		42445	=>	6544,
		42446	=>	6542,
		42447	=>	6540,
		42448	=>	6539,
		42449	=>	6537,
		42450	=>	6535,
		42451	=>	6533,
		42452	=>	6531,
		42453	=>	6529,
		42454	=>	6527,
		42455	=>	6525,
		42456	=>	6523,
		42457	=>	6522,
		42458	=>	6520,
		42459	=>	6518,
		42460	=>	6516,
		42461	=>	6514,
		42462	=>	6512,
		42463	=>	6510,
		42464	=>	6508,
		42465	=>	6507,
		42466	=>	6505,
		42467	=>	6503,
		42468	=>	6501,
		42469	=>	6499,
		42470	=>	6497,
		42471	=>	6495,
		42472	=>	6493,
		42473	=>	6492,
		42474	=>	6490,
		42475	=>	6488,
		42476	=>	6486,
		42477	=>	6484,
		42478	=>	6482,
		42479	=>	6480,
		42480	=>	6478,
		42481	=>	6476,
		42482	=>	6475,
		42483	=>	6473,
		42484	=>	6471,
		42485	=>	6469,
		42486	=>	6467,
		42487	=>	6465,
		42488	=>	6463,
		42489	=>	6462,
		42490	=>	6460,
		42491	=>	6458,
		42492	=>	6456,
		42493	=>	6454,
		42494	=>	6452,
		42495	=>	6450,
		42496	=>	6448,
		42497	=>	6447,
		42498	=>	6445,
		42499	=>	6443,
		42500	=>	6441,
		42501	=>	6439,
		42502	=>	6437,
		42503	=>	6435,
		42504	=>	6433,
		42505	=>	6432,
		42506	=>	6430,
		42507	=>	6428,
		42508	=>	6426,
		42509	=>	6424,
		42510	=>	6422,
		42511	=>	6420,
		42512	=>	6418,
		42513	=>	6417,
		42514	=>	6415,
		42515	=>	6413,
		42516	=>	6411,
		42517	=>	6409,
		42518	=>	6407,
		42519	=>	6405,
		42520	=>	6404,
		42521	=>	6402,
		42522	=>	6400,
		42523	=>	6398,
		42524	=>	6396,
		42525	=>	6394,
		42526	=>	6392,
		42527	=>	6390,
		42528	=>	6389,
		42529	=>	6387,
		42530	=>	6385,
		42531	=>	6383,
		42532	=>	6381,
		42533	=>	6379,
		42534	=>	6377,
		42535	=>	6376,
		42536	=>	6374,
		42537	=>	6372,
		42538	=>	6370,
		42539	=>	6368,
		42540	=>	6366,
		42541	=>	6364,
		42542	=>	6363,
		42543	=>	6361,
		42544	=>	6359,
		42545	=>	6357,
		42546	=>	6355,
		42547	=>	6353,
		42548	=>	6351,
		42549	=>	6350,
		42550	=>	6348,
		42551	=>	6346,
		42552	=>	6344,
		42553	=>	6342,
		42554	=>	6340,
		42555	=>	6338,
		42556	=>	6337,
		42557	=>	6335,
		42558	=>	6333,
		42559	=>	6331,
		42560	=>	6329,
		42561	=>	6327,
		42562	=>	6325,
		42563	=>	6324,
		42564	=>	6322,
		42565	=>	6320,
		42566	=>	6318,
		42567	=>	6316,
		42568	=>	6314,
		42569	=>	6312,
		42570	=>	6311,
		42571	=>	6309,
		42572	=>	6307,
		42573	=>	6305,
		42574	=>	6303,
		42575	=>	6301,
		42576	=>	6299,
		42577	=>	6298,
		42578	=>	6296,
		42579	=>	6294,
		42580	=>	6292,
		42581	=>	6290,
		42582	=>	6288,
		42583	=>	6287,
		42584	=>	6285,
		42585	=>	6283,
		42586	=>	6281,
		42587	=>	6279,
		42588	=>	6277,
		42589	=>	6275,
		42590	=>	6274,
		42591	=>	6272,
		42592	=>	6270,
		42593	=>	6268,
		42594	=>	6266,
		42595	=>	6264,
		42596	=>	6262,
		42597	=>	6261,
		42598	=>	6259,
		42599	=>	6257,
		42600	=>	6255,
		42601	=>	6253,
		42602	=>	6251,
		42603	=>	6250,
		42604	=>	6248,
		42605	=>	6246,
		42606	=>	6244,
		42607	=>	6242,
		42608	=>	6240,
		42609	=>	6238,
		42610	=>	6237,
		42611	=>	6235,
		42612	=>	6233,
		42613	=>	6231,
		42614	=>	6229,
		42615	=>	6227,
		42616	=>	6226,
		42617	=>	6224,
		42618	=>	6222,
		42619	=>	6220,
		42620	=>	6218,
		42621	=>	6216,
		42622	=>	6215,
		42623	=>	6213,
		42624	=>	6211,
		42625	=>	6209,
		42626	=>	6207,
		42627	=>	6205,
		42628	=>	6203,
		42629	=>	6202,
		42630	=>	6200,
		42631	=>	6198,
		42632	=>	6196,
		42633	=>	6194,
		42634	=>	6192,
		42635	=>	6191,
		42636	=>	6189,
		42637	=>	6187,
		42638	=>	6185,
		42639	=>	6183,
		42640	=>	6181,
		42641	=>	6180,
		42642	=>	6178,
		42643	=>	6176,
		42644	=>	6174,
		42645	=>	6172,
		42646	=>	6170,
		42647	=>	6169,
		42648	=>	6167,
		42649	=>	6165,
		42650	=>	6163,
		42651	=>	6161,
		42652	=>	6159,
		42653	=>	6158,
		42654	=>	6156,
		42655	=>	6154,
		42656	=>	6152,
		42657	=>	6150,
		42658	=>	6148,
		42659	=>	6147,
		42660	=>	6145,
		42661	=>	6143,
		42662	=>	6141,
		42663	=>	6139,
		42664	=>	6137,
		42665	=>	6136,
		42666	=>	6134,
		42667	=>	6132,
		42668	=>	6130,
		42669	=>	6128,
		42670	=>	6126,
		42671	=>	6125,
		42672	=>	6123,
		42673	=>	6121,
		42674	=>	6119,
		42675	=>	6117,
		42676	=>	6115,
		42677	=>	6114,
		42678	=>	6112,
		42679	=>	6110,
		42680	=>	6108,
		42681	=>	6106,
		42682	=>	6105,
		42683	=>	6103,
		42684	=>	6101,
		42685	=>	6099,
		42686	=>	6097,
		42687	=>	6095,
		42688	=>	6094,
		42689	=>	6092,
		42690	=>	6090,
		42691	=>	6088,
		42692	=>	6086,
		42693	=>	6084,
		42694	=>	6083,
		42695	=>	6081,
		42696	=>	6079,
		42697	=>	6077,
		42698	=>	6075,
		42699	=>	6074,
		42700	=>	6072,
		42701	=>	6070,
		42702	=>	6068,
		42703	=>	6066,
		42704	=>	6064,
		42705	=>	6063,
		42706	=>	6061,
		42707	=>	6059,
		42708	=>	6057,
		42709	=>	6055,
		42710	=>	6053,
		42711	=>	6052,
		42712	=>	6050,
		42713	=>	6048,
		42714	=>	6046,
		42715	=>	6044,
		42716	=>	6043,
		42717	=>	6041,
		42718	=>	6039,
		42719	=>	6037,
		42720	=>	6035,
		42721	=>	6033,
		42722	=>	6032,
		42723	=>	6030,
		42724	=>	6028,
		42725	=>	6026,
		42726	=>	6024,
		42727	=>	6023,
		42728	=>	6021,
		42729	=>	6019,
		42730	=>	6017,
		42731	=>	6015,
		42732	=>	6014,
		42733	=>	6012,
		42734	=>	6010,
		42735	=>	6008,
		42736	=>	6006,
		42737	=>	6004,
		42738	=>	6003,
		42739	=>	6001,
		42740	=>	5999,
		42741	=>	5997,
		42742	=>	5995,
		42743	=>	5994,
		42744	=>	5992,
		42745	=>	5990,
		42746	=>	5988,
		42747	=>	5986,
		42748	=>	5985,
		42749	=>	5983,
		42750	=>	5981,
		42751	=>	5979,
		42752	=>	5977,
		42753	=>	5975,
		42754	=>	5974,
		42755	=>	5972,
		42756	=>	5970,
		42757	=>	5968,
		42758	=>	5966,
		42759	=>	5965,
		42760	=>	5963,
		42761	=>	5961,
		42762	=>	5959,
		42763	=>	5957,
		42764	=>	5956,
		42765	=>	5954,
		42766	=>	5952,
		42767	=>	5950,
		42768	=>	5948,
		42769	=>	5947,
		42770	=>	5945,
		42771	=>	5943,
		42772	=>	5941,
		42773	=>	5939,
		42774	=>	5938,
		42775	=>	5936,
		42776	=>	5934,
		42777	=>	5932,
		42778	=>	5930,
		42779	=>	5929,
		42780	=>	5927,
		42781	=>	5925,
		42782	=>	5923,
		42783	=>	5921,
		42784	=>	5920,
		42785	=>	5918,
		42786	=>	5916,
		42787	=>	5914,
		42788	=>	5912,
		42789	=>	5911,
		42790	=>	5909,
		42791	=>	5907,
		42792	=>	5905,
		42793	=>	5903,
		42794	=>	5902,
		42795	=>	5900,
		42796	=>	5898,
		42797	=>	5896,
		42798	=>	5894,
		42799	=>	5893,
		42800	=>	5891,
		42801	=>	5889,
		42802	=>	5887,
		42803	=>	5885,
		42804	=>	5884,
		42805	=>	5882,
		42806	=>	5880,
		42807	=>	5878,
		42808	=>	5876,
		42809	=>	5875,
		42810	=>	5873,
		42811	=>	5871,
		42812	=>	5869,
		42813	=>	5867,
		42814	=>	5866,
		42815	=>	5864,
		42816	=>	5862,
		42817	=>	5860,
		42818	=>	5858,
		42819	=>	5857,
		42820	=>	5855,
		42821	=>	5853,
		42822	=>	5851,
		42823	=>	5849,
		42824	=>	5848,
		42825	=>	5846,
		42826	=>	5844,
		42827	=>	5842,
		42828	=>	5841,
		42829	=>	5839,
		42830	=>	5837,
		42831	=>	5835,
		42832	=>	5833,
		42833	=>	5832,
		42834	=>	5830,
		42835	=>	5828,
		42836	=>	5826,
		42837	=>	5824,
		42838	=>	5823,
		42839	=>	5821,
		42840	=>	5819,
		42841	=>	5817,
		42842	=>	5815,
		42843	=>	5814,
		42844	=>	5812,
		42845	=>	5810,
		42846	=>	5808,
		42847	=>	5807,
		42848	=>	5805,
		42849	=>	5803,
		42850	=>	5801,
		42851	=>	5799,
		42852	=>	5798,
		42853	=>	5796,
		42854	=>	5794,
		42855	=>	5792,
		42856	=>	5790,
		42857	=>	5789,
		42858	=>	5787,
		42859	=>	5785,
		42860	=>	5783,
		42861	=>	5782,
		42862	=>	5780,
		42863	=>	5778,
		42864	=>	5776,
		42865	=>	5774,
		42866	=>	5773,
		42867	=>	5771,
		42868	=>	5769,
		42869	=>	5767,
		42870	=>	5766,
		42871	=>	5764,
		42872	=>	5762,
		42873	=>	5760,
		42874	=>	5758,
		42875	=>	5757,
		42876	=>	5755,
		42877	=>	5753,
		42878	=>	5751,
		42879	=>	5750,
		42880	=>	5748,
		42881	=>	5746,
		42882	=>	5744,
		42883	=>	5742,
		42884	=>	5741,
		42885	=>	5739,
		42886	=>	5737,
		42887	=>	5735,
		42888	=>	5734,
		42889	=>	5732,
		42890	=>	5730,
		42891	=>	5728,
		42892	=>	5726,
		42893	=>	5725,
		42894	=>	5723,
		42895	=>	5721,
		42896	=>	5719,
		42897	=>	5718,
		42898	=>	5716,
		42899	=>	5714,
		42900	=>	5712,
		42901	=>	5711,
		42902	=>	5709,
		42903	=>	5707,
		42904	=>	5705,
		42905	=>	5703,
		42906	=>	5702,
		42907	=>	5700,
		42908	=>	5698,
		42909	=>	5696,
		42910	=>	5695,
		42911	=>	5693,
		42912	=>	5691,
		42913	=>	5689,
		42914	=>	5687,
		42915	=>	5686,
		42916	=>	5684,
		42917	=>	5682,
		42918	=>	5680,
		42919	=>	5679,
		42920	=>	5677,
		42921	=>	5675,
		42922	=>	5673,
		42923	=>	5672,
		42924	=>	5670,
		42925	=>	5668,
		42926	=>	5666,
		42927	=>	5665,
		42928	=>	5663,
		42929	=>	5661,
		42930	=>	5659,
		42931	=>	5657,
		42932	=>	5656,
		42933	=>	5654,
		42934	=>	5652,
		42935	=>	5650,
		42936	=>	5649,
		42937	=>	5647,
		42938	=>	5645,
		42939	=>	5643,
		42940	=>	5642,
		42941	=>	5640,
		42942	=>	5638,
		42943	=>	5636,
		42944	=>	5635,
		42945	=>	5633,
		42946	=>	5631,
		42947	=>	5629,
		42948	=>	5627,
		42949	=>	5626,
		42950	=>	5624,
		42951	=>	5622,
		42952	=>	5620,
		42953	=>	5619,
		42954	=>	5617,
		42955	=>	5615,
		42956	=>	5613,
		42957	=>	5612,
		42958	=>	5610,
		42959	=>	5608,
		42960	=>	5606,
		42961	=>	5605,
		42962	=>	5603,
		42963	=>	5601,
		42964	=>	5599,
		42965	=>	5598,
		42966	=>	5596,
		42967	=>	5594,
		42968	=>	5592,
		42969	=>	5591,
		42970	=>	5589,
		42971	=>	5587,
		42972	=>	5585,
		42973	=>	5584,
		42974	=>	5582,
		42975	=>	5580,
		42976	=>	5578,
		42977	=>	5577,
		42978	=>	5575,
		42979	=>	5573,
		42980	=>	5571,
		42981	=>	5570,
		42982	=>	5568,
		42983	=>	5566,
		42984	=>	5564,
		42985	=>	5563,
		42986	=>	5561,
		42987	=>	5559,
		42988	=>	5557,
		42989	=>	5556,
		42990	=>	5554,
		42991	=>	5552,
		42992	=>	5550,
		42993	=>	5549,
		42994	=>	5547,
		42995	=>	5545,
		42996	=>	5543,
		42997	=>	5542,
		42998	=>	5540,
		42999	=>	5538,
		43000	=>	5536,
		43001	=>	5535,
		43002	=>	5533,
		43003	=>	5531,
		43004	=>	5529,
		43005	=>	5528,
		43006	=>	5526,
		43007	=>	5524,
		43008	=>	5522,
		43009	=>	5521,
		43010	=>	5519,
		43011	=>	5517,
		43012	=>	5515,
		43013	=>	5514,
		43014	=>	5512,
		43015	=>	5510,
		43016	=>	5508,
		43017	=>	5507,
		43018	=>	5505,
		43019	=>	5503,
		43020	=>	5501,
		43021	=>	5500,
		43022	=>	5498,
		43023	=>	5496,
		43024	=>	5494,
		43025	=>	5493,
		43026	=>	5491,
		43027	=>	5489,
		43028	=>	5487,
		43029	=>	5486,
		43030	=>	5484,
		43031	=>	5482,
		43032	=>	5481,
		43033	=>	5479,
		43034	=>	5477,
		43035	=>	5475,
		43036	=>	5474,
		43037	=>	5472,
		43038	=>	5470,
		43039	=>	5468,
		43040	=>	5467,
		43041	=>	5465,
		43042	=>	5463,
		43043	=>	5461,
		43044	=>	5460,
		43045	=>	5458,
		43046	=>	5456,
		43047	=>	5454,
		43048	=>	5453,
		43049	=>	5451,
		43050	=>	5449,
		43051	=>	5448,
		43052	=>	5446,
		43053	=>	5444,
		43054	=>	5442,
		43055	=>	5441,
		43056	=>	5439,
		43057	=>	5437,
		43058	=>	5435,
		43059	=>	5434,
		43060	=>	5432,
		43061	=>	5430,
		43062	=>	5428,
		43063	=>	5427,
		43064	=>	5425,
		43065	=>	5423,
		43066	=>	5422,
		43067	=>	5420,
		43068	=>	5418,
		43069	=>	5416,
		43070	=>	5415,
		43071	=>	5413,
		43072	=>	5411,
		43073	=>	5409,
		43074	=>	5408,
		43075	=>	5406,
		43076	=>	5404,
		43077	=>	5402,
		43078	=>	5401,
		43079	=>	5399,
		43080	=>	5397,
		43081	=>	5396,
		43082	=>	5394,
		43083	=>	5392,
		43084	=>	5390,
		43085	=>	5389,
		43086	=>	5387,
		43087	=>	5385,
		43088	=>	5383,
		43089	=>	5382,
		43090	=>	5380,
		43091	=>	5378,
		43092	=>	5377,
		43093	=>	5375,
		43094	=>	5373,
		43095	=>	5371,
		43096	=>	5370,
		43097	=>	5368,
		43098	=>	5366,
		43099	=>	5365,
		43100	=>	5363,
		43101	=>	5361,
		43102	=>	5359,
		43103	=>	5358,
		43104	=>	5356,
		43105	=>	5354,
		43106	=>	5352,
		43107	=>	5351,
		43108	=>	5349,
		43109	=>	5347,
		43110	=>	5346,
		43111	=>	5344,
		43112	=>	5342,
		43113	=>	5340,
		43114	=>	5339,
		43115	=>	5337,
		43116	=>	5335,
		43117	=>	5334,
		43118	=>	5332,
		43119	=>	5330,
		43120	=>	5328,
		43121	=>	5327,
		43122	=>	5325,
		43123	=>	5323,
		43124	=>	5322,
		43125	=>	5320,
		43126	=>	5318,
		43127	=>	5316,
		43128	=>	5315,
		43129	=>	5313,
		43130	=>	5311,
		43131	=>	5310,
		43132	=>	5308,
		43133	=>	5306,
		43134	=>	5304,
		43135	=>	5303,
		43136	=>	5301,
		43137	=>	5299,
		43138	=>	5298,
		43139	=>	5296,
		43140	=>	5294,
		43141	=>	5292,
		43142	=>	5291,
		43143	=>	5289,
		43144	=>	5287,
		43145	=>	5286,
		43146	=>	5284,
		43147	=>	5282,
		43148	=>	5280,
		43149	=>	5279,
		43150	=>	5277,
		43151	=>	5275,
		43152	=>	5274,
		43153	=>	5272,
		43154	=>	5270,
		43155	=>	5268,
		43156	=>	5267,
		43157	=>	5265,
		43158	=>	5263,
		43159	=>	5262,
		43160	=>	5260,
		43161	=>	5258,
		43162	=>	5257,
		43163	=>	5255,
		43164	=>	5253,
		43165	=>	5251,
		43166	=>	5250,
		43167	=>	5248,
		43168	=>	5246,
		43169	=>	5245,
		43170	=>	5243,
		43171	=>	5241,
		43172	=>	5239,
		43173	=>	5238,
		43174	=>	5236,
		43175	=>	5234,
		43176	=>	5233,
		43177	=>	5231,
		43178	=>	5229,
		43179	=>	5228,
		43180	=>	5226,
		43181	=>	5224,
		43182	=>	5222,
		43183	=>	5221,
		43184	=>	5219,
		43185	=>	5217,
		43186	=>	5216,
		43187	=>	5214,
		43188	=>	5212,
		43189	=>	5211,
		43190	=>	5209,
		43191	=>	5207,
		43192	=>	5205,
		43193	=>	5204,
		43194	=>	5202,
		43195	=>	5200,
		43196	=>	5199,
		43197	=>	5197,
		43198	=>	5195,
		43199	=>	5194,
		43200	=>	5192,
		43201	=>	5190,
		43202	=>	5188,
		43203	=>	5187,
		43204	=>	5185,
		43205	=>	5183,
		43206	=>	5182,
		43207	=>	5180,
		43208	=>	5178,
		43209	=>	5177,
		43210	=>	5175,
		43211	=>	5173,
		43212	=>	5172,
		43213	=>	5170,
		43214	=>	5168,
		43215	=>	5166,
		43216	=>	5165,
		43217	=>	5163,
		43218	=>	5161,
		43219	=>	5160,
		43220	=>	5158,
		43221	=>	5156,
		43222	=>	5155,
		43223	=>	5153,
		43224	=>	5151,
		43225	=>	5150,
		43226	=>	5148,
		43227	=>	5146,
		43228	=>	5144,
		43229	=>	5143,
		43230	=>	5141,
		43231	=>	5139,
		43232	=>	5138,
		43233	=>	5136,
		43234	=>	5134,
		43235	=>	5133,
		43236	=>	5131,
		43237	=>	5129,
		43238	=>	5128,
		43239	=>	5126,
		43240	=>	5124,
		43241	=>	5122,
		43242	=>	5121,
		43243	=>	5119,
		43244	=>	5117,
		43245	=>	5116,
		43246	=>	5114,
		43247	=>	5112,
		43248	=>	5111,
		43249	=>	5109,
		43250	=>	5107,
		43251	=>	5106,
		43252	=>	5104,
		43253	=>	5102,
		43254	=>	5101,
		43255	=>	5099,
		43256	=>	5097,
		43257	=>	5096,
		43258	=>	5094,
		43259	=>	5092,
		43260	=>	5090,
		43261	=>	5089,
		43262	=>	5087,
		43263	=>	5085,
		43264	=>	5084,
		43265	=>	5082,
		43266	=>	5080,
		43267	=>	5079,
		43268	=>	5077,
		43269	=>	5075,
		43270	=>	5074,
		43271	=>	5072,
		43272	=>	5070,
		43273	=>	5069,
		43274	=>	5067,
		43275	=>	5065,
		43276	=>	5064,
		43277	=>	5062,
		43278	=>	5060,
		43279	=>	5059,
		43280	=>	5057,
		43281	=>	5055,
		43282	=>	5054,
		43283	=>	5052,
		43284	=>	5050,
		43285	=>	5049,
		43286	=>	5047,
		43287	=>	5045,
		43288	=>	5043,
		43289	=>	5042,
		43290	=>	5040,
		43291	=>	5038,
		43292	=>	5037,
		43293	=>	5035,
		43294	=>	5033,
		43295	=>	5032,
		43296	=>	5030,
		43297	=>	5028,
		43298	=>	5027,
		43299	=>	5025,
		43300	=>	5023,
		43301	=>	5022,
		43302	=>	5020,
		43303	=>	5018,
		43304	=>	5017,
		43305	=>	5015,
		43306	=>	5013,
		43307	=>	5012,
		43308	=>	5010,
		43309	=>	5008,
		43310	=>	5007,
		43311	=>	5005,
		43312	=>	5003,
		43313	=>	5002,
		43314	=>	5000,
		43315	=>	4998,
		43316	=>	4997,
		43317	=>	4995,
		43318	=>	4993,
		43319	=>	4992,
		43320	=>	4990,
		43321	=>	4988,
		43322	=>	4987,
		43323	=>	4985,
		43324	=>	4983,
		43325	=>	4982,
		43326	=>	4980,
		43327	=>	4978,
		43328	=>	4977,
		43329	=>	4975,
		43330	=>	4973,
		43331	=>	4972,
		43332	=>	4970,
		43333	=>	4968,
		43334	=>	4967,
		43335	=>	4965,
		43336	=>	4963,
		43337	=>	4962,
		43338	=>	4960,
		43339	=>	4958,
		43340	=>	4957,
		43341	=>	4955,
		43342	=>	4953,
		43343	=>	4952,
		43344	=>	4950,
		43345	=>	4948,
		43346	=>	4947,
		43347	=>	4945,
		43348	=>	4943,
		43349	=>	4942,
		43350	=>	4940,
		43351	=>	4939,
		43352	=>	4937,
		43353	=>	4935,
		43354	=>	4934,
		43355	=>	4932,
		43356	=>	4930,
		43357	=>	4929,
		43358	=>	4927,
		43359	=>	4925,
		43360	=>	4924,
		43361	=>	4922,
		43362	=>	4920,
		43363	=>	4919,
		43364	=>	4917,
		43365	=>	4915,
		43366	=>	4914,
		43367	=>	4912,
		43368	=>	4910,
		43369	=>	4909,
		43370	=>	4907,
		43371	=>	4905,
		43372	=>	4904,
		43373	=>	4902,
		43374	=>	4900,
		43375	=>	4899,
		43376	=>	4897,
		43377	=>	4895,
		43378	=>	4894,
		43379	=>	4892,
		43380	=>	4891,
		43381	=>	4889,
		43382	=>	4887,
		43383	=>	4886,
		43384	=>	4884,
		43385	=>	4882,
		43386	=>	4881,
		43387	=>	4879,
		43388	=>	4877,
		43389	=>	4876,
		43390	=>	4874,
		43391	=>	4872,
		43392	=>	4871,
		43393	=>	4869,
		43394	=>	4867,
		43395	=>	4866,
		43396	=>	4864,
		43397	=>	4862,
		43398	=>	4861,
		43399	=>	4859,
		43400	=>	4858,
		43401	=>	4856,
		43402	=>	4854,
		43403	=>	4853,
		43404	=>	4851,
		43405	=>	4849,
		43406	=>	4848,
		43407	=>	4846,
		43408	=>	4844,
		43409	=>	4843,
		43410	=>	4841,
		43411	=>	4839,
		43412	=>	4838,
		43413	=>	4836,
		43414	=>	4835,
		43415	=>	4833,
		43416	=>	4831,
		43417	=>	4830,
		43418	=>	4828,
		43419	=>	4826,
		43420	=>	4825,
		43421	=>	4823,
		43422	=>	4821,
		43423	=>	4820,
		43424	=>	4818,
		43425	=>	4816,
		43426	=>	4815,
		43427	=>	4813,
		43428	=>	4812,
		43429	=>	4810,
		43430	=>	4808,
		43431	=>	4807,
		43432	=>	4805,
		43433	=>	4803,
		43434	=>	4802,
		43435	=>	4800,
		43436	=>	4798,
		43437	=>	4797,
		43438	=>	4795,
		43439	=>	4794,
		43440	=>	4792,
		43441	=>	4790,
		43442	=>	4789,
		43443	=>	4787,
		43444	=>	4785,
		43445	=>	4784,
		43446	=>	4782,
		43447	=>	4780,
		43448	=>	4779,
		43449	=>	4777,
		43450	=>	4776,
		43451	=>	4774,
		43452	=>	4772,
		43453	=>	4771,
		43454	=>	4769,
		43455	=>	4767,
		43456	=>	4766,
		43457	=>	4764,
		43458	=>	4763,
		43459	=>	4761,
		43460	=>	4759,
		43461	=>	4758,
		43462	=>	4756,
		43463	=>	4754,
		43464	=>	4753,
		43465	=>	4751,
		43466	=>	4749,
		43467	=>	4748,
		43468	=>	4746,
		43469	=>	4745,
		43470	=>	4743,
		43471	=>	4741,
		43472	=>	4740,
		43473	=>	4738,
		43474	=>	4736,
		43475	=>	4735,
		43476	=>	4733,
		43477	=>	4732,
		43478	=>	4730,
		43479	=>	4728,
		43480	=>	4727,
		43481	=>	4725,
		43482	=>	4723,
		43483	=>	4722,
		43484	=>	4720,
		43485	=>	4719,
		43486	=>	4717,
		43487	=>	4715,
		43488	=>	4714,
		43489	=>	4712,
		43490	=>	4710,
		43491	=>	4709,
		43492	=>	4707,
		43493	=>	4706,
		43494	=>	4704,
		43495	=>	4702,
		43496	=>	4701,
		43497	=>	4699,
		43498	=>	4697,
		43499	=>	4696,
		43500	=>	4694,
		43501	=>	4693,
		43502	=>	4691,
		43503	=>	4689,
		43504	=>	4688,
		43505	=>	4686,
		43506	=>	4685,
		43507	=>	4683,
		43508	=>	4681,
		43509	=>	4680,
		43510	=>	4678,
		43511	=>	4676,
		43512	=>	4675,
		43513	=>	4673,
		43514	=>	4672,
		43515	=>	4670,
		43516	=>	4668,
		43517	=>	4667,
		43518	=>	4665,
		43519	=>	4663,
		43520	=>	4662,
		43521	=>	4660,
		43522	=>	4659,
		43523	=>	4657,
		43524	=>	4655,
		43525	=>	4654,
		43526	=>	4652,
		43527	=>	4651,
		43528	=>	4649,
		43529	=>	4647,
		43530	=>	4646,
		43531	=>	4644,
		43532	=>	4643,
		43533	=>	4641,
		43534	=>	4639,
		43535	=>	4638,
		43536	=>	4636,
		43537	=>	4634,
		43538	=>	4633,
		43539	=>	4631,
		43540	=>	4630,
		43541	=>	4628,
		43542	=>	4626,
		43543	=>	4625,
		43544	=>	4623,
		43545	=>	4622,
		43546	=>	4620,
		43547	=>	4618,
		43548	=>	4617,
		43549	=>	4615,
		43550	=>	4614,
		43551	=>	4612,
		43552	=>	4610,
		43553	=>	4609,
		43554	=>	4607,
		43555	=>	4606,
		43556	=>	4604,
		43557	=>	4602,
		43558	=>	4601,
		43559	=>	4599,
		43560	=>	4597,
		43561	=>	4596,
		43562	=>	4594,
		43563	=>	4593,
		43564	=>	4591,
		43565	=>	4589,
		43566	=>	4588,
		43567	=>	4586,
		43568	=>	4585,
		43569	=>	4583,
		43570	=>	4581,
		43571	=>	4580,
		43572	=>	4578,
		43573	=>	4577,
		43574	=>	4575,
		43575	=>	4573,
		43576	=>	4572,
		43577	=>	4570,
		43578	=>	4569,
		43579	=>	4567,
		43580	=>	4565,
		43581	=>	4564,
		43582	=>	4562,
		43583	=>	4561,
		43584	=>	4559,
		43585	=>	4557,
		43586	=>	4556,
		43587	=>	4554,
		43588	=>	4553,
		43589	=>	4551,
		43590	=>	4549,
		43591	=>	4548,
		43592	=>	4546,
		43593	=>	4545,
		43594	=>	4543,
		43595	=>	4541,
		43596	=>	4540,
		43597	=>	4538,
		43598	=>	4537,
		43599	=>	4535,
		43600	=>	4533,
		43601	=>	4532,
		43602	=>	4530,
		43603	=>	4529,
		43604	=>	4527,
		43605	=>	4526,
		43606	=>	4524,
		43607	=>	4522,
		43608	=>	4521,
		43609	=>	4519,
		43610	=>	4518,
		43611	=>	4516,
		43612	=>	4514,
		43613	=>	4513,
		43614	=>	4511,
		43615	=>	4510,
		43616	=>	4508,
		43617	=>	4506,
		43618	=>	4505,
		43619	=>	4503,
		43620	=>	4502,
		43621	=>	4500,
		43622	=>	4498,
		43623	=>	4497,
		43624	=>	4495,
		43625	=>	4494,
		43626	=>	4492,
		43627	=>	4491,
		43628	=>	4489,
		43629	=>	4487,
		43630	=>	4486,
		43631	=>	4484,
		43632	=>	4483,
		43633	=>	4481,
		43634	=>	4479,
		43635	=>	4478,
		43636	=>	4476,
		43637	=>	4475,
		43638	=>	4473,
		43639	=>	4472,
		43640	=>	4470,
		43641	=>	4468,
		43642	=>	4467,
		43643	=>	4465,
		43644	=>	4464,
		43645	=>	4462,
		43646	=>	4460,
		43647	=>	4459,
		43648	=>	4457,
		43649	=>	4456,
		43650	=>	4454,
		43651	=>	4453,
		43652	=>	4451,
		43653	=>	4449,
		43654	=>	4448,
		43655	=>	4446,
		43656	=>	4445,
		43657	=>	4443,
		43658	=>	4441,
		43659	=>	4440,
		43660	=>	4438,
		43661	=>	4437,
		43662	=>	4435,
		43663	=>	4434,
		43664	=>	4432,
		43665	=>	4430,
		43666	=>	4429,
		43667	=>	4427,
		43668	=>	4426,
		43669	=>	4424,
		43670	=>	4423,
		43671	=>	4421,
		43672	=>	4419,
		43673	=>	4418,
		43674	=>	4416,
		43675	=>	4415,
		43676	=>	4413,
		43677	=>	4412,
		43678	=>	4410,
		43679	=>	4408,
		43680	=>	4407,
		43681	=>	4405,
		43682	=>	4404,
		43683	=>	4402,
		43684	=>	4400,
		43685	=>	4399,
		43686	=>	4397,
		43687	=>	4396,
		43688	=>	4394,
		43689	=>	4393,
		43690	=>	4391,
		43691	=>	4389,
		43692	=>	4388,
		43693	=>	4386,
		43694	=>	4385,
		43695	=>	4383,
		43696	=>	4382,
		43697	=>	4380,
		43698	=>	4379,
		43699	=>	4377,
		43700	=>	4375,
		43701	=>	4374,
		43702	=>	4372,
		43703	=>	4371,
		43704	=>	4369,
		43705	=>	4368,
		43706	=>	4366,
		43707	=>	4364,
		43708	=>	4363,
		43709	=>	4361,
		43710	=>	4360,
		43711	=>	4358,
		43712	=>	4357,
		43713	=>	4355,
		43714	=>	4353,
		43715	=>	4352,
		43716	=>	4350,
		43717	=>	4349,
		43718	=>	4347,
		43719	=>	4346,
		43720	=>	4344,
		43721	=>	4342,
		43722	=>	4341,
		43723	=>	4339,
		43724	=>	4338,
		43725	=>	4336,
		43726	=>	4335,
		43727	=>	4333,
		43728	=>	4332,
		43729	=>	4330,
		43730	=>	4328,
		43731	=>	4327,
		43732	=>	4325,
		43733	=>	4324,
		43734	=>	4322,
		43735	=>	4321,
		43736	=>	4319,
		43737	=>	4318,
		43738	=>	4316,
		43739	=>	4314,
		43740	=>	4313,
		43741	=>	4311,
		43742	=>	4310,
		43743	=>	4308,
		43744	=>	4307,
		43745	=>	4305,
		43746	=>	4303,
		43747	=>	4302,
		43748	=>	4300,
		43749	=>	4299,
		43750	=>	4297,
		43751	=>	4296,
		43752	=>	4294,
		43753	=>	4293,
		43754	=>	4291,
		43755	=>	4289,
		43756	=>	4288,
		43757	=>	4286,
		43758	=>	4285,
		43759	=>	4283,
		43760	=>	4282,
		43761	=>	4280,
		43762	=>	4279,
		43763	=>	4277,
		43764	=>	4276,
		43765	=>	4274,
		43766	=>	4272,
		43767	=>	4271,
		43768	=>	4269,
		43769	=>	4268,
		43770	=>	4266,
		43771	=>	4265,
		43772	=>	4263,
		43773	=>	4262,
		43774	=>	4260,
		43775	=>	4258,
		43776	=>	4257,
		43777	=>	4255,
		43778	=>	4254,
		43779	=>	4252,
		43780	=>	4251,
		43781	=>	4249,
		43782	=>	4248,
		43783	=>	4246,
		43784	=>	4245,
		43785	=>	4243,
		43786	=>	4241,
		43787	=>	4240,
		43788	=>	4238,
		43789	=>	4237,
		43790	=>	4235,
		43791	=>	4234,
		43792	=>	4232,
		43793	=>	4231,
		43794	=>	4229,
		43795	=>	4228,
		43796	=>	4226,
		43797	=>	4224,
		43798	=>	4223,
		43799	=>	4221,
		43800	=>	4220,
		43801	=>	4218,
		43802	=>	4217,
		43803	=>	4215,
		43804	=>	4214,
		43805	=>	4212,
		43806	=>	4211,
		43807	=>	4209,
		43808	=>	4208,
		43809	=>	4206,
		43810	=>	4204,
		43811	=>	4203,
		43812	=>	4201,
		43813	=>	4200,
		43814	=>	4198,
		43815	=>	4197,
		43816	=>	4195,
		43817	=>	4194,
		43818	=>	4192,
		43819	=>	4191,
		43820	=>	4189,
		43821	=>	4188,
		43822	=>	4186,
		43823	=>	4184,
		43824	=>	4183,
		43825	=>	4181,
		43826	=>	4180,
		43827	=>	4178,
		43828	=>	4177,
		43829	=>	4175,
		43830	=>	4174,
		43831	=>	4172,
		43832	=>	4171,
		43833	=>	4169,
		43834	=>	4168,
		43835	=>	4166,
		43836	=>	4164,
		43837	=>	4163,
		43838	=>	4161,
		43839	=>	4160,
		43840	=>	4158,
		43841	=>	4157,
		43842	=>	4155,
		43843	=>	4154,
		43844	=>	4152,
		43845	=>	4151,
		43846	=>	4149,
		43847	=>	4148,
		43848	=>	4146,
		43849	=>	4145,
		43850	=>	4143,
		43851	=>	4142,
		43852	=>	4140,
		43853	=>	4138,
		43854	=>	4137,
		43855	=>	4135,
		43856	=>	4134,
		43857	=>	4132,
		43858	=>	4131,
		43859	=>	4129,
		43860	=>	4128,
		43861	=>	4126,
		43862	=>	4125,
		43863	=>	4123,
		43864	=>	4122,
		43865	=>	4120,
		43866	=>	4119,
		43867	=>	4117,
		43868	=>	4116,
		43869	=>	4114,
		43870	=>	4113,
		43871	=>	4111,
		43872	=>	4109,
		43873	=>	4108,
		43874	=>	4106,
		43875	=>	4105,
		43876	=>	4103,
		43877	=>	4102,
		43878	=>	4100,
		43879	=>	4099,
		43880	=>	4097,
		43881	=>	4096,
		43882	=>	4094,
		43883	=>	4093,
		43884	=>	4091,
		43885	=>	4090,
		43886	=>	4088,
		43887	=>	4087,
		43888	=>	4085,
		43889	=>	4084,
		43890	=>	4082,
		43891	=>	4081,
		43892	=>	4079,
		43893	=>	4078,
		43894	=>	4076,
		43895	=>	4075,
		43896	=>	4073,
		43897	=>	4071,
		43898	=>	4070,
		43899	=>	4068,
		43900	=>	4067,
		43901	=>	4065,
		43902	=>	4064,
		43903	=>	4062,
		43904	=>	4061,
		43905	=>	4059,
		43906	=>	4058,
		43907	=>	4056,
		43908	=>	4055,
		43909	=>	4053,
		43910	=>	4052,
		43911	=>	4050,
		43912	=>	4049,
		43913	=>	4047,
		43914	=>	4046,
		43915	=>	4044,
		43916	=>	4043,
		43917	=>	4041,
		43918	=>	4040,
		43919	=>	4038,
		43920	=>	4037,
		43921	=>	4035,
		43922	=>	4034,
		43923	=>	4032,
		43924	=>	4031,
		43925	=>	4029,
		43926	=>	4028,
		43927	=>	4026,
		43928	=>	4025,
		43929	=>	4023,
		43930	=>	4022,
		43931	=>	4020,
		43932	=>	4019,
		43933	=>	4017,
		43934	=>	4016,
		43935	=>	4014,
		43936	=>	4013,
		43937	=>	4011,
		43938	=>	4010,
		43939	=>	4008,
		43940	=>	4007,
		43941	=>	4005,
		43942	=>	4004,
		43943	=>	4002,
		43944	=>	4000,
		43945	=>	3999,
		43946	=>	3997,
		43947	=>	3996,
		43948	=>	3994,
		43949	=>	3993,
		43950	=>	3991,
		43951	=>	3990,
		43952	=>	3988,
		43953	=>	3987,
		43954	=>	3985,
		43955	=>	3984,
		43956	=>	3982,
		43957	=>	3981,
		43958	=>	3979,
		43959	=>	3978,
		43960	=>	3976,
		43961	=>	3975,
		43962	=>	3973,
		43963	=>	3972,
		43964	=>	3970,
		43965	=>	3969,
		43966	=>	3967,
		43967	=>	3966,
		43968	=>	3964,
		43969	=>	3963,
		43970	=>	3961,
		43971	=>	3960,
		43972	=>	3958,
		43973	=>	3957,
		43974	=>	3955,
		43975	=>	3954,
		43976	=>	3952,
		43977	=>	3951,
		43978	=>	3950,
		43979	=>	3948,
		43980	=>	3947,
		43981	=>	3945,
		43982	=>	3944,
		43983	=>	3942,
		43984	=>	3941,
		43985	=>	3939,
		43986	=>	3938,
		43987	=>	3936,
		43988	=>	3935,
		43989	=>	3933,
		43990	=>	3932,
		43991	=>	3930,
		43992	=>	3929,
		43993	=>	3927,
		43994	=>	3926,
		43995	=>	3924,
		43996	=>	3923,
		43997	=>	3921,
		43998	=>	3920,
		43999	=>	3918,
		44000	=>	3917,
		44001	=>	3915,
		44002	=>	3914,
		44003	=>	3912,
		44004	=>	3911,
		44005	=>	3909,
		44006	=>	3908,
		44007	=>	3906,
		44008	=>	3905,
		44009	=>	3903,
		44010	=>	3902,
		44011	=>	3900,
		44012	=>	3899,
		44013	=>	3897,
		44014	=>	3896,
		44015	=>	3894,
		44016	=>	3893,
		44017	=>	3891,
		44018	=>	3890,
		44019	=>	3888,
		44020	=>	3887,
		44021	=>	3885,
		44022	=>	3884,
		44023	=>	3882,
		44024	=>	3881,
		44025	=>	3880,
		44026	=>	3878,
		44027	=>	3877,
		44028	=>	3875,
		44029	=>	3874,
		44030	=>	3872,
		44031	=>	3871,
		44032	=>	3869,
		44033	=>	3868,
		44034	=>	3866,
		44035	=>	3865,
		44036	=>	3863,
		44037	=>	3862,
		44038	=>	3860,
		44039	=>	3859,
		44040	=>	3857,
		44041	=>	3856,
		44042	=>	3854,
		44043	=>	3853,
		44044	=>	3851,
		44045	=>	3850,
		44046	=>	3848,
		44047	=>	3847,
		44048	=>	3845,
		44049	=>	3844,
		44050	=>	3843,
		44051	=>	3841,
		44052	=>	3840,
		44053	=>	3838,
		44054	=>	3837,
		44055	=>	3835,
		44056	=>	3834,
		44057	=>	3832,
		44058	=>	3831,
		44059	=>	3829,
		44060	=>	3828,
		44061	=>	3826,
		44062	=>	3825,
		44063	=>	3823,
		44064	=>	3822,
		44065	=>	3820,
		44066	=>	3819,
		44067	=>	3817,
		44068	=>	3816,
		44069	=>	3815,
		44070	=>	3813,
		44071	=>	3812,
		44072	=>	3810,
		44073	=>	3809,
		44074	=>	3807,
		44075	=>	3806,
		44076	=>	3804,
		44077	=>	3803,
		44078	=>	3801,
		44079	=>	3800,
		44080	=>	3798,
		44081	=>	3797,
		44082	=>	3795,
		44083	=>	3794,
		44084	=>	3792,
		44085	=>	3791,
		44086	=>	3790,
		44087	=>	3788,
		44088	=>	3787,
		44089	=>	3785,
		44090	=>	3784,
		44091	=>	3782,
		44092	=>	3781,
		44093	=>	3779,
		44094	=>	3778,
		44095	=>	3776,
		44096	=>	3775,
		44097	=>	3773,
		44098	=>	3772,
		44099	=>	3771,
		44100	=>	3769,
		44101	=>	3768,
		44102	=>	3766,
		44103	=>	3765,
		44104	=>	3763,
		44105	=>	3762,
		44106	=>	3760,
		44107	=>	3759,
		44108	=>	3757,
		44109	=>	3756,
		44110	=>	3754,
		44111	=>	3753,
		44112	=>	3752,
		44113	=>	3750,
		44114	=>	3749,
		44115	=>	3747,
		44116	=>	3746,
		44117	=>	3744,
		44118	=>	3743,
		44119	=>	3741,
		44120	=>	3740,
		44121	=>	3738,
		44122	=>	3737,
		44123	=>	3735,
		44124	=>	3734,
		44125	=>	3733,
		44126	=>	3731,
		44127	=>	3730,
		44128	=>	3728,
		44129	=>	3727,
		44130	=>	3725,
		44131	=>	3724,
		44132	=>	3722,
		44133	=>	3721,
		44134	=>	3719,
		44135	=>	3718,
		44136	=>	3717,
		44137	=>	3715,
		44138	=>	3714,
		44139	=>	3712,
		44140	=>	3711,
		44141	=>	3709,
		44142	=>	3708,
		44143	=>	3706,
		44144	=>	3705,
		44145	=>	3704,
		44146	=>	3702,
		44147	=>	3701,
		44148	=>	3699,
		44149	=>	3698,
		44150	=>	3696,
		44151	=>	3695,
		44152	=>	3693,
		44153	=>	3692,
		44154	=>	3690,
		44155	=>	3689,
		44156	=>	3688,
		44157	=>	3686,
		44158	=>	3685,
		44159	=>	3683,
		44160	=>	3682,
		44161	=>	3680,
		44162	=>	3679,
		44163	=>	3677,
		44164	=>	3676,
		44165	=>	3675,
		44166	=>	3673,
		44167	=>	3672,
		44168	=>	3670,
		44169	=>	3669,
		44170	=>	3667,
		44171	=>	3666,
		44172	=>	3664,
		44173	=>	3663,
		44174	=>	3662,
		44175	=>	3660,
		44176	=>	3659,
		44177	=>	3657,
		44178	=>	3656,
		44179	=>	3654,
		44180	=>	3653,
		44181	=>	3651,
		44182	=>	3650,
		44183	=>	3649,
		44184	=>	3647,
		44185	=>	3646,
		44186	=>	3644,
		44187	=>	3643,
		44188	=>	3641,
		44189	=>	3640,
		44190	=>	3638,
		44191	=>	3637,
		44192	=>	3636,
		44193	=>	3634,
		44194	=>	3633,
		44195	=>	3631,
		44196	=>	3630,
		44197	=>	3628,
		44198	=>	3627,
		44199	=>	3626,
		44200	=>	3624,
		44201	=>	3623,
		44202	=>	3621,
		44203	=>	3620,
		44204	=>	3618,
		44205	=>	3617,
		44206	=>	3615,
		44207	=>	3614,
		44208	=>	3613,
		44209	=>	3611,
		44210	=>	3610,
		44211	=>	3608,
		44212	=>	3607,
		44213	=>	3605,
		44214	=>	3604,
		44215	=>	3603,
		44216	=>	3601,
		44217	=>	3600,
		44218	=>	3598,
		44219	=>	3597,
		44220	=>	3595,
		44221	=>	3594,
		44222	=>	3593,
		44223	=>	3591,
		44224	=>	3590,
		44225	=>	3588,
		44226	=>	3587,
		44227	=>	3585,
		44228	=>	3584,
		44229	=>	3583,
		44230	=>	3581,
		44231	=>	3580,
		44232	=>	3578,
		44233	=>	3577,
		44234	=>	3575,
		44235	=>	3574,
		44236	=>	3573,
		44237	=>	3571,
		44238	=>	3570,
		44239	=>	3568,
		44240	=>	3567,
		44241	=>	3565,
		44242	=>	3564,
		44243	=>	3563,
		44244	=>	3561,
		44245	=>	3560,
		44246	=>	3558,
		44247	=>	3557,
		44248	=>	3555,
		44249	=>	3554,
		44250	=>	3553,
		44251	=>	3551,
		44252	=>	3550,
		44253	=>	3548,
		44254	=>	3547,
		44255	=>	3546,
		44256	=>	3544,
		44257	=>	3543,
		44258	=>	3541,
		44259	=>	3540,
		44260	=>	3538,
		44261	=>	3537,
		44262	=>	3536,
		44263	=>	3534,
		44264	=>	3533,
		44265	=>	3531,
		44266	=>	3530,
		44267	=>	3528,
		44268	=>	3527,
		44269	=>	3526,
		44270	=>	3524,
		44271	=>	3523,
		44272	=>	3521,
		44273	=>	3520,
		44274	=>	3519,
		44275	=>	3517,
		44276	=>	3516,
		44277	=>	3514,
		44278	=>	3513,
		44279	=>	3511,
		44280	=>	3510,
		44281	=>	3509,
		44282	=>	3507,
		44283	=>	3506,
		44284	=>	3504,
		44285	=>	3503,
		44286	=>	3502,
		44287	=>	3500,
		44288	=>	3499,
		44289	=>	3497,
		44290	=>	3496,
		44291	=>	3495,
		44292	=>	3493,
		44293	=>	3492,
		44294	=>	3490,
		44295	=>	3489,
		44296	=>	3487,
		44297	=>	3486,
		44298	=>	3485,
		44299	=>	3483,
		44300	=>	3482,
		44301	=>	3480,
		44302	=>	3479,
		44303	=>	3478,
		44304	=>	3476,
		44305	=>	3475,
		44306	=>	3473,
		44307	=>	3472,
		44308	=>	3471,
		44309	=>	3469,
		44310	=>	3468,
		44311	=>	3466,
		44312	=>	3465,
		44313	=>	3464,
		44314	=>	3462,
		44315	=>	3461,
		44316	=>	3459,
		44317	=>	3458,
		44318	=>	3457,
		44319	=>	3455,
		44320	=>	3454,
		44321	=>	3452,
		44322	=>	3451,
		44323	=>	3450,
		44324	=>	3448,
		44325	=>	3447,
		44326	=>	3445,
		44327	=>	3444,
		44328	=>	3442,
		44329	=>	3441,
		44330	=>	3440,
		44331	=>	3438,
		44332	=>	3437,
		44333	=>	3435,
		44334	=>	3434,
		44335	=>	3433,
		44336	=>	3431,
		44337	=>	3430,
		44338	=>	3428,
		44339	=>	3427,
		44340	=>	3426,
		44341	=>	3424,
		44342	=>	3423,
		44343	=>	3421,
		44344	=>	3420,
		44345	=>	3419,
		44346	=>	3417,
		44347	=>	3416,
		44348	=>	3415,
		44349	=>	3413,
		44350	=>	3412,
		44351	=>	3410,
		44352	=>	3409,
		44353	=>	3408,
		44354	=>	3406,
		44355	=>	3405,
		44356	=>	3403,
		44357	=>	3402,
		44358	=>	3401,
		44359	=>	3399,
		44360	=>	3398,
		44361	=>	3396,
		44362	=>	3395,
		44363	=>	3394,
		44364	=>	3392,
		44365	=>	3391,
		44366	=>	3389,
		44367	=>	3388,
		44368	=>	3387,
		44369	=>	3385,
		44370	=>	3384,
		44371	=>	3382,
		44372	=>	3381,
		44373	=>	3380,
		44374	=>	3378,
		44375	=>	3377,
		44376	=>	3376,
		44377	=>	3374,
		44378	=>	3373,
		44379	=>	3371,
		44380	=>	3370,
		44381	=>	3369,
		44382	=>	3367,
		44383	=>	3366,
		44384	=>	3364,
		44385	=>	3363,
		44386	=>	3362,
		44387	=>	3360,
		44388	=>	3359,
		44389	=>	3357,
		44390	=>	3356,
		44391	=>	3355,
		44392	=>	3353,
		44393	=>	3352,
		44394	=>	3351,
		44395	=>	3349,
		44396	=>	3348,
		44397	=>	3346,
		44398	=>	3345,
		44399	=>	3344,
		44400	=>	3342,
		44401	=>	3341,
		44402	=>	3340,
		44403	=>	3338,
		44404	=>	3337,
		44405	=>	3335,
		44406	=>	3334,
		44407	=>	3333,
		44408	=>	3331,
		44409	=>	3330,
		44410	=>	3328,
		44411	=>	3327,
		44412	=>	3326,
		44413	=>	3324,
		44414	=>	3323,
		44415	=>	3322,
		44416	=>	3320,
		44417	=>	3319,
		44418	=>	3317,
		44419	=>	3316,
		44420	=>	3315,
		44421	=>	3313,
		44422	=>	3312,
		44423	=>	3311,
		44424	=>	3309,
		44425	=>	3308,
		44426	=>	3306,
		44427	=>	3305,
		44428	=>	3304,
		44429	=>	3302,
		44430	=>	3301,
		44431	=>	3300,
		44432	=>	3298,
		44433	=>	3297,
		44434	=>	3295,
		44435	=>	3294,
		44436	=>	3293,
		44437	=>	3291,
		44438	=>	3290,
		44439	=>	3289,
		44440	=>	3287,
		44441	=>	3286,
		44442	=>	3284,
		44443	=>	3283,
		44444	=>	3282,
		44445	=>	3280,
		44446	=>	3279,
		44447	=>	3278,
		44448	=>	3276,
		44449	=>	3275,
		44450	=>	3273,
		44451	=>	3272,
		44452	=>	3271,
		44453	=>	3269,
		44454	=>	3268,
		44455	=>	3267,
		44456	=>	3265,
		44457	=>	3264,
		44458	=>	3263,
		44459	=>	3261,
		44460	=>	3260,
		44461	=>	3258,
		44462	=>	3257,
		44463	=>	3256,
		44464	=>	3254,
		44465	=>	3253,
		44466	=>	3252,
		44467	=>	3250,
		44468	=>	3249,
		44469	=>	3248,
		44470	=>	3246,
		44471	=>	3245,
		44472	=>	3243,
		44473	=>	3242,
		44474	=>	3241,
		44475	=>	3239,
		44476	=>	3238,
		44477	=>	3237,
		44478	=>	3235,
		44479	=>	3234,
		44480	=>	3233,
		44481	=>	3231,
		44482	=>	3230,
		44483	=>	3228,
		44484	=>	3227,
		44485	=>	3226,
		44486	=>	3224,
		44487	=>	3223,
		44488	=>	3222,
		44489	=>	3220,
		44490	=>	3219,
		44491	=>	3218,
		44492	=>	3216,
		44493	=>	3215,
		44494	=>	3214,
		44495	=>	3212,
		44496	=>	3211,
		44497	=>	3209,
		44498	=>	3208,
		44499	=>	3207,
		44500	=>	3205,
		44501	=>	3204,
		44502	=>	3203,
		44503	=>	3201,
		44504	=>	3200,
		44505	=>	3199,
		44506	=>	3197,
		44507	=>	3196,
		44508	=>	3195,
		44509	=>	3193,
		44510	=>	3192,
		44511	=>	3191,
		44512	=>	3189,
		44513	=>	3188,
		44514	=>	3186,
		44515	=>	3185,
		44516	=>	3184,
		44517	=>	3182,
		44518	=>	3181,
		44519	=>	3180,
		44520	=>	3178,
		44521	=>	3177,
		44522	=>	3176,
		44523	=>	3174,
		44524	=>	3173,
		44525	=>	3172,
		44526	=>	3170,
		44527	=>	3169,
		44528	=>	3168,
		44529	=>	3166,
		44530	=>	3165,
		44531	=>	3164,
		44532	=>	3162,
		44533	=>	3161,
		44534	=>	3159,
		44535	=>	3158,
		44536	=>	3157,
		44537	=>	3155,
		44538	=>	3154,
		44539	=>	3153,
		44540	=>	3151,
		44541	=>	3150,
		44542	=>	3149,
		44543	=>	3147,
		44544	=>	3146,
		44545	=>	3145,
		44546	=>	3143,
		44547	=>	3142,
		44548	=>	3141,
		44549	=>	3139,
		44550	=>	3138,
		44551	=>	3137,
		44552	=>	3135,
		44553	=>	3134,
		44554	=>	3133,
		44555	=>	3131,
		44556	=>	3130,
		44557	=>	3129,
		44558	=>	3127,
		44559	=>	3126,
		44560	=>	3125,
		44561	=>	3123,
		44562	=>	3122,
		44563	=>	3121,
		44564	=>	3119,
		44565	=>	3118,
		44566	=>	3117,
		44567	=>	3115,
		44568	=>	3114,
		44569	=>	3113,
		44570	=>	3111,
		44571	=>	3110,
		44572	=>	3109,
		44573	=>	3107,
		44574	=>	3106,
		44575	=>	3105,
		44576	=>	3103,
		44577	=>	3102,
		44578	=>	3101,
		44579	=>	3099,
		44580	=>	3098,
		44581	=>	3097,
		44582	=>	3095,
		44583	=>	3094,
		44584	=>	3093,
		44585	=>	3091,
		44586	=>	3090,
		44587	=>	3089,
		44588	=>	3087,
		44589	=>	3086,
		44590	=>	3085,
		44591	=>	3083,
		44592	=>	3082,
		44593	=>	3081,
		44594	=>	3079,
		44595	=>	3078,
		44596	=>	3077,
		44597	=>	3075,
		44598	=>	3074,
		44599	=>	3073,
		44600	=>	3071,
		44601	=>	3070,
		44602	=>	3069,
		44603	=>	3067,
		44604	=>	3066,
		44605	=>	3065,
		44606	=>	3063,
		44607	=>	3062,
		44608	=>	3061,
		44609	=>	3059,
		44610	=>	3058,
		44611	=>	3057,
		44612	=>	3055,
		44613	=>	3054,
		44614	=>	3053,
		44615	=>	3051,
		44616	=>	3050,
		44617	=>	3049,
		44618	=>	3047,
		44619	=>	3046,
		44620	=>	3045,
		44621	=>	3043,
		44622	=>	3042,
		44623	=>	3041,
		44624	=>	3039,
		44625	=>	3038,
		44626	=>	3037,
		44627	=>	3035,
		44628	=>	3034,
		44629	=>	3033,
		44630	=>	3032,
		44631	=>	3030,
		44632	=>	3029,
		44633	=>	3028,
		44634	=>	3026,
		44635	=>	3025,
		44636	=>	3024,
		44637	=>	3022,
		44638	=>	3021,
		44639	=>	3020,
		44640	=>	3018,
		44641	=>	3017,
		44642	=>	3016,
		44643	=>	3014,
		44644	=>	3013,
		44645	=>	3012,
		44646	=>	3010,
		44647	=>	3009,
		44648	=>	3008,
		44649	=>	3006,
		44650	=>	3005,
		44651	=>	3004,
		44652	=>	3003,
		44653	=>	3001,
		44654	=>	3000,
		44655	=>	2999,
		44656	=>	2997,
		44657	=>	2996,
		44658	=>	2995,
		44659	=>	2993,
		44660	=>	2992,
		44661	=>	2991,
		44662	=>	2989,
		44663	=>	2988,
		44664	=>	2987,
		44665	=>	2986,
		44666	=>	2984,
		44667	=>	2983,
		44668	=>	2982,
		44669	=>	2980,
		44670	=>	2979,
		44671	=>	2978,
		44672	=>	2976,
		44673	=>	2975,
		44674	=>	2974,
		44675	=>	2972,
		44676	=>	2971,
		44677	=>	2970,
		44678	=>	2968,
		44679	=>	2967,
		44680	=>	2966,
		44681	=>	2965,
		44682	=>	2963,
		44683	=>	2962,
		44684	=>	2961,
		44685	=>	2959,
		44686	=>	2958,
		44687	=>	2957,
		44688	=>	2955,
		44689	=>	2954,
		44690	=>	2953,
		44691	=>	2952,
		44692	=>	2950,
		44693	=>	2949,
		44694	=>	2948,
		44695	=>	2946,
		44696	=>	2945,
		44697	=>	2944,
		44698	=>	2942,
		44699	=>	2941,
		44700	=>	2940,
		44701	=>	2939,
		44702	=>	2937,
		44703	=>	2936,
		44704	=>	2935,
		44705	=>	2933,
		44706	=>	2932,
		44707	=>	2931,
		44708	=>	2929,
		44709	=>	2928,
		44710	=>	2927,
		44711	=>	2926,
		44712	=>	2924,
		44713	=>	2923,
		44714	=>	2922,
		44715	=>	2920,
		44716	=>	2919,
		44717	=>	2918,
		44718	=>	2916,
		44719	=>	2915,
		44720	=>	2914,
		44721	=>	2913,
		44722	=>	2911,
		44723	=>	2910,
		44724	=>	2909,
		44725	=>	2907,
		44726	=>	2906,
		44727	=>	2905,
		44728	=>	2904,
		44729	=>	2902,
		44730	=>	2901,
		44731	=>	2900,
		44732	=>	2898,
		44733	=>	2897,
		44734	=>	2896,
		44735	=>	2894,
		44736	=>	2893,
		44737	=>	2892,
		44738	=>	2891,
		44739	=>	2889,
		44740	=>	2888,
		44741	=>	2887,
		44742	=>	2885,
		44743	=>	2884,
		44744	=>	2883,
		44745	=>	2882,
		44746	=>	2880,
		44747	=>	2879,
		44748	=>	2878,
		44749	=>	2876,
		44750	=>	2875,
		44751	=>	2874,
		44752	=>	2873,
		44753	=>	2871,
		44754	=>	2870,
		44755	=>	2869,
		44756	=>	2867,
		44757	=>	2866,
		44758	=>	2865,
		44759	=>	2864,
		44760	=>	2862,
		44761	=>	2861,
		44762	=>	2860,
		44763	=>	2858,
		44764	=>	2857,
		44765	=>	2856,
		44766	=>	2855,
		44767	=>	2853,
		44768	=>	2852,
		44769	=>	2851,
		44770	=>	2849,
		44771	=>	2848,
		44772	=>	2847,
		44773	=>	2846,
		44774	=>	2844,
		44775	=>	2843,
		44776	=>	2842,
		44777	=>	2840,
		44778	=>	2839,
		44779	=>	2838,
		44780	=>	2837,
		44781	=>	2835,
		44782	=>	2834,
		44783	=>	2833,
		44784	=>	2832,
		44785	=>	2830,
		44786	=>	2829,
		44787	=>	2828,
		44788	=>	2826,
		44789	=>	2825,
		44790	=>	2824,
		44791	=>	2823,
		44792	=>	2821,
		44793	=>	2820,
		44794	=>	2819,
		44795	=>	2818,
		44796	=>	2816,
		44797	=>	2815,
		44798	=>	2814,
		44799	=>	2812,
		44800	=>	2811,
		44801	=>	2810,
		44802	=>	2809,
		44803	=>	2807,
		44804	=>	2806,
		44805	=>	2805,
		44806	=>	2803,
		44807	=>	2802,
		44808	=>	2801,
		44809	=>	2800,
		44810	=>	2798,
		44811	=>	2797,
		44812	=>	2796,
		44813	=>	2795,
		44814	=>	2793,
		44815	=>	2792,
		44816	=>	2791,
		44817	=>	2790,
		44818	=>	2788,
		44819	=>	2787,
		44820	=>	2786,
		44821	=>	2784,
		44822	=>	2783,
		44823	=>	2782,
		44824	=>	2781,
		44825	=>	2779,
		44826	=>	2778,
		44827	=>	2777,
		44828	=>	2776,
		44829	=>	2774,
		44830	=>	2773,
		44831	=>	2772,
		44832	=>	2771,
		44833	=>	2769,
		44834	=>	2768,
		44835	=>	2767,
		44836	=>	2765,
		44837	=>	2764,
		44838	=>	2763,
		44839	=>	2762,
		44840	=>	2760,
		44841	=>	2759,
		44842	=>	2758,
		44843	=>	2757,
		44844	=>	2755,
		44845	=>	2754,
		44846	=>	2753,
		44847	=>	2752,
		44848	=>	2750,
		44849	=>	2749,
		44850	=>	2748,
		44851	=>	2747,
		44852	=>	2745,
		44853	=>	2744,
		44854	=>	2743,
		44855	=>	2742,
		44856	=>	2740,
		44857	=>	2739,
		44858	=>	2738,
		44859	=>	2736,
		44860	=>	2735,
		44861	=>	2734,
		44862	=>	2733,
		44863	=>	2731,
		44864	=>	2730,
		44865	=>	2729,
		44866	=>	2728,
		44867	=>	2726,
		44868	=>	2725,
		44869	=>	2724,
		44870	=>	2723,
		44871	=>	2721,
		44872	=>	2720,
		44873	=>	2719,
		44874	=>	2718,
		44875	=>	2716,
		44876	=>	2715,
		44877	=>	2714,
		44878	=>	2713,
		44879	=>	2711,
		44880	=>	2710,
		44881	=>	2709,
		44882	=>	2708,
		44883	=>	2706,
		44884	=>	2705,
		44885	=>	2704,
		44886	=>	2703,
		44887	=>	2701,
		44888	=>	2700,
		44889	=>	2699,
		44890	=>	2698,
		44891	=>	2696,
		44892	=>	2695,
		44893	=>	2694,
		44894	=>	2693,
		44895	=>	2691,
		44896	=>	2690,
		44897	=>	2689,
		44898	=>	2688,
		44899	=>	2686,
		44900	=>	2685,
		44901	=>	2684,
		44902	=>	2683,
		44903	=>	2681,
		44904	=>	2680,
		44905	=>	2679,
		44906	=>	2678,
		44907	=>	2676,
		44908	=>	2675,
		44909	=>	2674,
		44910	=>	2673,
		44911	=>	2672,
		44912	=>	2670,
		44913	=>	2669,
		44914	=>	2668,
		44915	=>	2667,
		44916	=>	2665,
		44917	=>	2664,
		44918	=>	2663,
		44919	=>	2662,
		44920	=>	2660,
		44921	=>	2659,
		44922	=>	2658,
		44923	=>	2657,
		44924	=>	2655,
		44925	=>	2654,
		44926	=>	2653,
		44927	=>	2652,
		44928	=>	2650,
		44929	=>	2649,
		44930	=>	2648,
		44931	=>	2647,
		44932	=>	2645,
		44933	=>	2644,
		44934	=>	2643,
		44935	=>	2642,
		44936	=>	2641,
		44937	=>	2639,
		44938	=>	2638,
		44939	=>	2637,
		44940	=>	2636,
		44941	=>	2634,
		44942	=>	2633,
		44943	=>	2632,
		44944	=>	2631,
		44945	=>	2629,
		44946	=>	2628,
		44947	=>	2627,
		44948	=>	2626,
		44949	=>	2625,
		44950	=>	2623,
		44951	=>	2622,
		44952	=>	2621,
		44953	=>	2620,
		44954	=>	2618,
		44955	=>	2617,
		44956	=>	2616,
		44957	=>	2615,
		44958	=>	2613,
		44959	=>	2612,
		44960	=>	2611,
		44961	=>	2610,
		44962	=>	2609,
		44963	=>	2607,
		44964	=>	2606,
		44965	=>	2605,
		44966	=>	2604,
		44967	=>	2602,
		44968	=>	2601,
		44969	=>	2600,
		44970	=>	2599,
		44971	=>	2597,
		44972	=>	2596,
		44973	=>	2595,
		44974	=>	2594,
		44975	=>	2593,
		44976	=>	2591,
		44977	=>	2590,
		44978	=>	2589,
		44979	=>	2588,
		44980	=>	2586,
		44981	=>	2585,
		44982	=>	2584,
		44983	=>	2583,
		44984	=>	2582,
		44985	=>	2580,
		44986	=>	2579,
		44987	=>	2578,
		44988	=>	2577,
		44989	=>	2575,
		44990	=>	2574,
		44991	=>	2573,
		44992	=>	2572,
		44993	=>	2571,
		44994	=>	2569,
		44995	=>	2568,
		44996	=>	2567,
		44997	=>	2566,
		44998	=>	2564,
		44999	=>	2563,
		45000	=>	2562,
		45001	=>	2561,
		45002	=>	2560,
		45003	=>	2558,
		45004	=>	2557,
		45005	=>	2556,
		45006	=>	2555,
		45007	=>	2554,
		45008	=>	2552,
		45009	=>	2551,
		45010	=>	2550,
		45011	=>	2549,
		45012	=>	2547,
		45013	=>	2546,
		45014	=>	2545,
		45015	=>	2544,
		45016	=>	2543,
		45017	=>	2541,
		45018	=>	2540,
		45019	=>	2539,
		45020	=>	2538,
		45021	=>	2537,
		45022	=>	2535,
		45023	=>	2534,
		45024	=>	2533,
		45025	=>	2532,
		45026	=>	2530,
		45027	=>	2529,
		45028	=>	2528,
		45029	=>	2527,
		45030	=>	2526,
		45031	=>	2524,
		45032	=>	2523,
		45033	=>	2522,
		45034	=>	2521,
		45035	=>	2520,
		45036	=>	2518,
		45037	=>	2517,
		45038	=>	2516,
		45039	=>	2515,
		45040	=>	2514,
		45041	=>	2512,
		45042	=>	2511,
		45043	=>	2510,
		45044	=>	2509,
		45045	=>	2508,
		45046	=>	2506,
		45047	=>	2505,
		45048	=>	2504,
		45049	=>	2503,
		45050	=>	2501,
		45051	=>	2500,
		45052	=>	2499,
		45053	=>	2498,
		45054	=>	2497,
		45055	=>	2495,
		45056	=>	2494,
		45057	=>	2493,
		45058	=>	2492,
		45059	=>	2491,
		45060	=>	2489,
		45061	=>	2488,
		45062	=>	2487,
		45063	=>	2486,
		45064	=>	2485,
		45065	=>	2483,
		45066	=>	2482,
		45067	=>	2481,
		45068	=>	2480,
		45069	=>	2479,
		45070	=>	2477,
		45071	=>	2476,
		45072	=>	2475,
		45073	=>	2474,
		45074	=>	2473,
		45075	=>	2471,
		45076	=>	2470,
		45077	=>	2469,
		45078	=>	2468,
		45079	=>	2467,
		45080	=>	2466,
		45081	=>	2464,
		45082	=>	2463,
		45083	=>	2462,
		45084	=>	2461,
		45085	=>	2460,
		45086	=>	2458,
		45087	=>	2457,
		45088	=>	2456,
		45089	=>	2455,
		45090	=>	2454,
		45091	=>	2452,
		45092	=>	2451,
		45093	=>	2450,
		45094	=>	2449,
		45095	=>	2448,
		45096	=>	2446,
		45097	=>	2445,
		45098	=>	2444,
		45099	=>	2443,
		45100	=>	2442,
		45101	=>	2440,
		45102	=>	2439,
		45103	=>	2438,
		45104	=>	2437,
		45105	=>	2436,
		45106	=>	2435,
		45107	=>	2433,
		45108	=>	2432,
		45109	=>	2431,
		45110	=>	2430,
		45111	=>	2429,
		45112	=>	2427,
		45113	=>	2426,
		45114	=>	2425,
		45115	=>	2424,
		45116	=>	2423,
		45117	=>	2421,
		45118	=>	2420,
		45119	=>	2419,
		45120	=>	2418,
		45121	=>	2417,
		45122	=>	2416,
		45123	=>	2414,
		45124	=>	2413,
		45125	=>	2412,
		45126	=>	2411,
		45127	=>	2410,
		45128	=>	2408,
		45129	=>	2407,
		45130	=>	2406,
		45131	=>	2405,
		45132	=>	2404,
		45133	=>	2403,
		45134	=>	2401,
		45135	=>	2400,
		45136	=>	2399,
		45137	=>	2398,
		45138	=>	2397,
		45139	=>	2395,
		45140	=>	2394,
		45141	=>	2393,
		45142	=>	2392,
		45143	=>	2391,
		45144	=>	2390,
		45145	=>	2388,
		45146	=>	2387,
		45147	=>	2386,
		45148	=>	2385,
		45149	=>	2384,
		45150	=>	2382,
		45151	=>	2381,
		45152	=>	2380,
		45153	=>	2379,
		45154	=>	2378,
		45155	=>	2377,
		45156	=>	2375,
		45157	=>	2374,
		45158	=>	2373,
		45159	=>	2372,
		45160	=>	2371,
		45161	=>	2370,
		45162	=>	2368,
		45163	=>	2367,
		45164	=>	2366,
		45165	=>	2365,
		45166	=>	2364,
		45167	=>	2363,
		45168	=>	2361,
		45169	=>	2360,
		45170	=>	2359,
		45171	=>	2358,
		45172	=>	2357,
		45173	=>	2356,
		45174	=>	2354,
		45175	=>	2353,
		45176	=>	2352,
		45177	=>	2351,
		45178	=>	2350,
		45179	=>	2349,
		45180	=>	2347,
		45181	=>	2346,
		45182	=>	2345,
		45183	=>	2344,
		45184	=>	2343,
		45185	=>	2342,
		45186	=>	2340,
		45187	=>	2339,
		45188	=>	2338,
		45189	=>	2337,
		45190	=>	2336,
		45191	=>	2335,
		45192	=>	2333,
		45193	=>	2332,
		45194	=>	2331,
		45195	=>	2330,
		45196	=>	2329,
		45197	=>	2328,
		45198	=>	2326,
		45199	=>	2325,
		45200	=>	2324,
		45201	=>	2323,
		45202	=>	2322,
		45203	=>	2321,
		45204	=>	2319,
		45205	=>	2318,
		45206	=>	2317,
		45207	=>	2316,
		45208	=>	2315,
		45209	=>	2314,
		45210	=>	2312,
		45211	=>	2311,
		45212	=>	2310,
		45213	=>	2309,
		45214	=>	2308,
		45215	=>	2307,
		45216	=>	2305,
		45217	=>	2304,
		45218	=>	2303,
		45219	=>	2302,
		45220	=>	2301,
		45221	=>	2300,
		45222	=>	2299,
		45223	=>	2297,
		45224	=>	2296,
		45225	=>	2295,
		45226	=>	2294,
		45227	=>	2293,
		45228	=>	2292,
		45229	=>	2290,
		45230	=>	2289,
		45231	=>	2288,
		45232	=>	2287,
		45233	=>	2286,
		45234	=>	2285,
		45235	=>	2284,
		45236	=>	2282,
		45237	=>	2281,
		45238	=>	2280,
		45239	=>	2279,
		45240	=>	2278,
		45241	=>	2277,
		45242	=>	2275,
		45243	=>	2274,
		45244	=>	2273,
		45245	=>	2272,
		45246	=>	2271,
		45247	=>	2270,
		45248	=>	2269,
		45249	=>	2267,
		45250	=>	2266,
		45251	=>	2265,
		45252	=>	2264,
		45253	=>	2263,
		45254	=>	2262,
		45255	=>	2261,
		45256	=>	2259,
		45257	=>	2258,
		45258	=>	2257,
		45259	=>	2256,
		45260	=>	2255,
		45261	=>	2254,
		45262	=>	2253,
		45263	=>	2251,
		45264	=>	2250,
		45265	=>	2249,
		45266	=>	2248,
		45267	=>	2247,
		45268	=>	2246,
		45269	=>	2245,
		45270	=>	2243,
		45271	=>	2242,
		45272	=>	2241,
		45273	=>	2240,
		45274	=>	2239,
		45275	=>	2238,
		45276	=>	2237,
		45277	=>	2235,
		45278	=>	2234,
		45279	=>	2233,
		45280	=>	2232,
		45281	=>	2231,
		45282	=>	2230,
		45283	=>	2229,
		45284	=>	2227,
		45285	=>	2226,
		45286	=>	2225,
		45287	=>	2224,
		45288	=>	2223,
		45289	=>	2222,
		45290	=>	2221,
		45291	=>	2219,
		45292	=>	2218,
		45293	=>	2217,
		45294	=>	2216,
		45295	=>	2215,
		45296	=>	2214,
		45297	=>	2213,
		45298	=>	2212,
		45299	=>	2210,
		45300	=>	2209,
		45301	=>	2208,
		45302	=>	2207,
		45303	=>	2206,
		45304	=>	2205,
		45305	=>	2204,
		45306	=>	2202,
		45307	=>	2201,
		45308	=>	2200,
		45309	=>	2199,
		45310	=>	2198,
		45311	=>	2197,
		45312	=>	2196,
		45313	=>	2195,
		45314	=>	2193,
		45315	=>	2192,
		45316	=>	2191,
		45317	=>	2190,
		45318	=>	2189,
		45319	=>	2188,
		45320	=>	2187,
		45321	=>	2185,
		45322	=>	2184,
		45323	=>	2183,
		45324	=>	2182,
		45325	=>	2181,
		45326	=>	2180,
		45327	=>	2179,
		45328	=>	2178,
		45329	=>	2176,
		45330	=>	2175,
		45331	=>	2174,
		45332	=>	2173,
		45333	=>	2172,
		45334	=>	2171,
		45335	=>	2170,
		45336	=>	2169,
		45337	=>	2167,
		45338	=>	2166,
		45339	=>	2165,
		45340	=>	2164,
		45341	=>	2163,
		45342	=>	2162,
		45343	=>	2161,
		45344	=>	2160,
		45345	=>	2159,
		45346	=>	2157,
		45347	=>	2156,
		45348	=>	2155,
		45349	=>	2154,
		45350	=>	2153,
		45351	=>	2152,
		45352	=>	2151,
		45353	=>	2150,
		45354	=>	2148,
		45355	=>	2147,
		45356	=>	2146,
		45357	=>	2145,
		45358	=>	2144,
		45359	=>	2143,
		45360	=>	2142,
		45361	=>	2141,
		45362	=>	2139,
		45363	=>	2138,
		45364	=>	2137,
		45365	=>	2136,
		45366	=>	2135,
		45367	=>	2134,
		45368	=>	2133,
		45369	=>	2132,
		45370	=>	2131,
		45371	=>	2129,
		45372	=>	2128,
		45373	=>	2127,
		45374	=>	2126,
		45375	=>	2125,
		45376	=>	2124,
		45377	=>	2123,
		45378	=>	2122,
		45379	=>	2121,
		45380	=>	2119,
		45381	=>	2118,
		45382	=>	2117,
		45383	=>	2116,
		45384	=>	2115,
		45385	=>	2114,
		45386	=>	2113,
		45387	=>	2112,
		45388	=>	2111,
		45389	=>	2109,
		45390	=>	2108,
		45391	=>	2107,
		45392	=>	2106,
		45393	=>	2105,
		45394	=>	2104,
		45395	=>	2103,
		45396	=>	2102,
		45397	=>	2101,
		45398	=>	2099,
		45399	=>	2098,
		45400	=>	2097,
		45401	=>	2096,
		45402	=>	2095,
		45403	=>	2094,
		45404	=>	2093,
		45405	=>	2092,
		45406	=>	2091,
		45407	=>	2090,
		45408	=>	2088,
		45409	=>	2087,
		45410	=>	2086,
		45411	=>	2085,
		45412	=>	2084,
		45413	=>	2083,
		45414	=>	2082,
		45415	=>	2081,
		45416	=>	2080,
		45417	=>	2078,
		45418	=>	2077,
		45419	=>	2076,
		45420	=>	2075,
		45421	=>	2074,
		45422	=>	2073,
		45423	=>	2072,
		45424	=>	2071,
		45425	=>	2070,
		45426	=>	2069,
		45427	=>	2067,
		45428	=>	2066,
		45429	=>	2065,
		45430	=>	2064,
		45431	=>	2063,
		45432	=>	2062,
		45433	=>	2061,
		45434	=>	2060,
		45435	=>	2059,
		45436	=>	2058,
		45437	=>	2057,
		45438	=>	2055,
		45439	=>	2054,
		45440	=>	2053,
		45441	=>	2052,
		45442	=>	2051,
		45443	=>	2050,
		45444	=>	2049,
		45445	=>	2048,
		45446	=>	2047,
		45447	=>	2046,
		45448	=>	2044,
		45449	=>	2043,
		45450	=>	2042,
		45451	=>	2041,
		45452	=>	2040,
		45453	=>	2039,
		45454	=>	2038,
		45455	=>	2037,
		45456	=>	2036,
		45457	=>	2035,
		45458	=>	2034,
		45459	=>	2032,
		45460	=>	2031,
		45461	=>	2030,
		45462	=>	2029,
		45463	=>	2028,
		45464	=>	2027,
		45465	=>	2026,
		45466	=>	2025,
		45467	=>	2024,
		45468	=>	2023,
		45469	=>	2022,
		45470	=>	2021,
		45471	=>	2019,
		45472	=>	2018,
		45473	=>	2017,
		45474	=>	2016,
		45475	=>	2015,
		45476	=>	2014,
		45477	=>	2013,
		45478	=>	2012,
		45479	=>	2011,
		45480	=>	2010,
		45481	=>	2009,
		45482	=>	2008,
		45483	=>	2006,
		45484	=>	2005,
		45485	=>	2004,
		45486	=>	2003,
		45487	=>	2002,
		45488	=>	2001,
		45489	=>	2000,
		45490	=>	1999,
		45491	=>	1998,
		45492	=>	1997,
		45493	=>	1996,
		45494	=>	1995,
		45495	=>	1993,
		45496	=>	1992,
		45497	=>	1991,
		45498	=>	1990,
		45499	=>	1989,
		45500	=>	1988,
		45501	=>	1987,
		45502	=>	1986,
		45503	=>	1985,
		45504	=>	1984,
		45505	=>	1983,
		45506	=>	1982,
		45507	=>	1981,
		45508	=>	1979,
		45509	=>	1978,
		45510	=>	1977,
		45511	=>	1976,
		45512	=>	1975,
		45513	=>	1974,
		45514	=>	1973,
		45515	=>	1972,
		45516	=>	1971,
		45517	=>	1970,
		45518	=>	1969,
		45519	=>	1968,
		45520	=>	1967,
		45521	=>	1966,
		45522	=>	1964,
		45523	=>	1963,
		45524	=>	1962,
		45525	=>	1961,
		45526	=>	1960,
		45527	=>	1959,
		45528	=>	1958,
		45529	=>	1957,
		45530	=>	1956,
		45531	=>	1955,
		45532	=>	1954,
		45533	=>	1953,
		45534	=>	1952,
		45535	=>	1951,
		45536	=>	1949,
		45537	=>	1948,
		45538	=>	1947,
		45539	=>	1946,
		45540	=>	1945,
		45541	=>	1944,
		45542	=>	1943,
		45543	=>	1942,
		45544	=>	1941,
		45545	=>	1940,
		45546	=>	1939,
		45547	=>	1938,
		45548	=>	1937,
		45549	=>	1936,
		45550	=>	1935,
		45551	=>	1933,
		45552	=>	1932,
		45553	=>	1931,
		45554	=>	1930,
		45555	=>	1929,
		45556	=>	1928,
		45557	=>	1927,
		45558	=>	1926,
		45559	=>	1925,
		45560	=>	1924,
		45561	=>	1923,
		45562	=>	1922,
		45563	=>	1921,
		45564	=>	1920,
		45565	=>	1919,
		45566	=>	1918,
		45567	=>	1917,
		45568	=>	1915,
		45569	=>	1914,
		45570	=>	1913,
		45571	=>	1912,
		45572	=>	1911,
		45573	=>	1910,
		45574	=>	1909,
		45575	=>	1908,
		45576	=>	1907,
		45577	=>	1906,
		45578	=>	1905,
		45579	=>	1904,
		45580	=>	1903,
		45581	=>	1902,
		45582	=>	1901,
		45583	=>	1900,
		45584	=>	1899,
		45585	=>	1898,
		45586	=>	1896,
		45587	=>	1895,
		45588	=>	1894,
		45589	=>	1893,
		45590	=>	1892,
		45591	=>	1891,
		45592	=>	1890,
		45593	=>	1889,
		45594	=>	1888,
		45595	=>	1887,
		45596	=>	1886,
		45597	=>	1885,
		45598	=>	1884,
		45599	=>	1883,
		45600	=>	1882,
		45601	=>	1881,
		45602	=>	1880,
		45603	=>	1879,
		45604	=>	1878,
		45605	=>	1876,
		45606	=>	1875,
		45607	=>	1874,
		45608	=>	1873,
		45609	=>	1872,
		45610	=>	1871,
		45611	=>	1870,
		45612	=>	1869,
		45613	=>	1868,
		45614	=>	1867,
		45615	=>	1866,
		45616	=>	1865,
		45617	=>	1864,
		45618	=>	1863,
		45619	=>	1862,
		45620	=>	1861,
		45621	=>	1860,
		45622	=>	1859,
		45623	=>	1858,
		45624	=>	1857,
		45625	=>	1856,
		45626	=>	1855,
		45627	=>	1854,
		45628	=>	1852,
		45629	=>	1851,
		45630	=>	1850,
		45631	=>	1849,
		45632	=>	1848,
		45633	=>	1847,
		45634	=>	1846,
		45635	=>	1845,
		45636	=>	1844,
		45637	=>	1843,
		45638	=>	1842,
		45639	=>	1841,
		45640	=>	1840,
		45641	=>	1839,
		45642	=>	1838,
		45643	=>	1837,
		45644	=>	1836,
		45645	=>	1835,
		45646	=>	1834,
		45647	=>	1833,
		45648	=>	1832,
		45649	=>	1831,
		45650	=>	1830,
		45651	=>	1829,
		45652	=>	1828,
		45653	=>	1827,
		45654	=>	1825,
		45655	=>	1824,
		45656	=>	1823,
		45657	=>	1822,
		45658	=>	1821,
		45659	=>	1820,
		45660	=>	1819,
		45661	=>	1818,
		45662	=>	1817,
		45663	=>	1816,
		45664	=>	1815,
		45665	=>	1814,
		45666	=>	1813,
		45667	=>	1812,
		45668	=>	1811,
		45669	=>	1810,
		45670	=>	1809,
		45671	=>	1808,
		45672	=>	1807,
		45673	=>	1806,
		45674	=>	1805,
		45675	=>	1804,
		45676	=>	1803,
		45677	=>	1802,
		45678	=>	1801,
		45679	=>	1800,
		45680	=>	1799,
		45681	=>	1798,
		45682	=>	1797,
		45683	=>	1796,
		45684	=>	1795,
		45685	=>	1794,
		45686	=>	1793,
		45687	=>	1792,
		45688	=>	1790,
		45689	=>	1789,
		45690	=>	1788,
		45691	=>	1787,
		45692	=>	1786,
		45693	=>	1785,
		45694	=>	1784,
		45695	=>	1783,
		45696	=>	1782,
		45697	=>	1781,
		45698	=>	1780,
		45699	=>	1779,
		45700	=>	1778,
		45701	=>	1777,
		45702	=>	1776,
		45703	=>	1775,
		45704	=>	1774,
		45705	=>	1773,
		45706	=>	1772,
		45707	=>	1771,
		45708	=>	1770,
		45709	=>	1769,
		45710	=>	1768,
		45711	=>	1767,
		45712	=>	1766,
		45713	=>	1765,
		45714	=>	1764,
		45715	=>	1763,
		45716	=>	1762,
		45717	=>	1761,
		45718	=>	1760,
		45719	=>	1759,
		45720	=>	1758,
		45721	=>	1757,
		45722	=>	1756,
		45723	=>	1755,
		45724	=>	1754,
		45725	=>	1753,
		45726	=>	1752,
		45727	=>	1751,
		45728	=>	1750,
		45729	=>	1749,
		45730	=>	1748,
		45731	=>	1747,
		45732	=>	1746,
		45733	=>	1745,
		45734	=>	1744,
		45735	=>	1743,
		45736	=>	1742,
		45737	=>	1741,
		45738	=>	1740,
		45739	=>	1739,
		45740	=>	1738,
		45741	=>	1737,
		45742	=>	1736,
		45743	=>	1735,
		45744	=>	1734,
		45745	=>	1733,
		45746	=>	1732,
		45747	=>	1731,
		45748	=>	1730,
		45749	=>	1729,
		45750	=>	1728,
		45751	=>	1727,
		45752	=>	1726,
		45753	=>	1725,
		45754	=>	1724,
		45755	=>	1723,
		45756	=>	1722,
		45757	=>	1721,
		45758	=>	1719,
		45759	=>	1718,
		45760	=>	1717,
		45761	=>	1716,
		45762	=>	1715,
		45763	=>	1714,
		45764	=>	1713,
		45765	=>	1712,
		45766	=>	1711,
		45767	=>	1710,
		45768	=>	1709,
		45769	=>	1708,
		45770	=>	1707,
		45771	=>	1706,
		45772	=>	1705,
		45773	=>	1704,
		45774	=>	1703,
		45775	=>	1702,
		45776	=>	1701,
		45777	=>	1700,
		45778	=>	1699,
		45779	=>	1698,
		45780	=>	1697,
		45781	=>	1696,
		45782	=>	1695,
		45783	=>	1694,
		45784	=>	1693,
		45785	=>	1692,
		45786	=>	1691,
		45787	=>	1690,
		45788	=>	1689,
		45789	=>	1689,
		45790	=>	1688,
		45791	=>	1687,
		45792	=>	1686,
		45793	=>	1685,
		45794	=>	1684,
		45795	=>	1683,
		45796	=>	1682,
		45797	=>	1681,
		45798	=>	1680,
		45799	=>	1679,
		45800	=>	1678,
		45801	=>	1677,
		45802	=>	1676,
		45803	=>	1675,
		45804	=>	1674,
		45805	=>	1673,
		45806	=>	1672,
		45807	=>	1671,
		45808	=>	1670,
		45809	=>	1669,
		45810	=>	1668,
		45811	=>	1667,
		45812	=>	1666,
		45813	=>	1665,
		45814	=>	1664,
		45815	=>	1663,
		45816	=>	1662,
		45817	=>	1661,
		45818	=>	1660,
		45819	=>	1659,
		45820	=>	1658,
		45821	=>	1657,
		45822	=>	1656,
		45823	=>	1655,
		45824	=>	1654,
		45825	=>	1653,
		45826	=>	1652,
		45827	=>	1651,
		45828	=>	1650,
		45829	=>	1649,
		45830	=>	1648,
		45831	=>	1647,
		45832	=>	1646,
		45833	=>	1645,
		45834	=>	1644,
		45835	=>	1643,
		45836	=>	1642,
		45837	=>	1641,
		45838	=>	1640,
		45839	=>	1639,
		45840	=>	1638,
		45841	=>	1637,
		45842	=>	1636,
		45843	=>	1635,
		45844	=>	1634,
		45845	=>	1633,
		45846	=>	1632,
		45847	=>	1631,
		45848	=>	1630,
		45849	=>	1629,
		45850	=>	1628,
		45851	=>	1627,
		45852	=>	1626,
		45853	=>	1625,
		45854	=>	1624,
		45855	=>	1623,
		45856	=>	1622,
		45857	=>	1621,
		45858	=>	1620,
		45859	=>	1620,
		45860	=>	1619,
		45861	=>	1618,
		45862	=>	1617,
		45863	=>	1616,
		45864	=>	1615,
		45865	=>	1614,
		45866	=>	1613,
		45867	=>	1612,
		45868	=>	1611,
		45869	=>	1610,
		45870	=>	1609,
		45871	=>	1608,
		45872	=>	1607,
		45873	=>	1606,
		45874	=>	1605,
		45875	=>	1604,
		45876	=>	1603,
		45877	=>	1602,
		45878	=>	1601,
		45879	=>	1600,
		45880	=>	1599,
		45881	=>	1598,
		45882	=>	1597,
		45883	=>	1596,
		45884	=>	1595,
		45885	=>	1594,
		45886	=>	1593,
		45887	=>	1592,
		45888	=>	1591,
		45889	=>	1590,
		45890	=>	1589,
		45891	=>	1588,
		45892	=>	1587,
		45893	=>	1587,
		45894	=>	1586,
		45895	=>	1585,
		45896	=>	1584,
		45897	=>	1583,
		45898	=>	1582,
		45899	=>	1581,
		45900	=>	1580,
		45901	=>	1579,
		45902	=>	1578,
		45903	=>	1577,
		45904	=>	1576,
		45905	=>	1575,
		45906	=>	1574,
		45907	=>	1573,
		45908	=>	1572,
		45909	=>	1571,
		45910	=>	1570,
		45911	=>	1569,
		45912	=>	1568,
		45913	=>	1567,
		45914	=>	1566,
		45915	=>	1565,
		45916	=>	1564,
		45917	=>	1563,
		45918	=>	1562,
		45919	=>	1562,
		45920	=>	1561,
		45921	=>	1560,
		45922	=>	1559,
		45923	=>	1558,
		45924	=>	1557,
		45925	=>	1556,
		45926	=>	1555,
		45927	=>	1554,
		45928	=>	1553,
		45929	=>	1552,
		45930	=>	1551,
		45931	=>	1550,
		45932	=>	1549,
		45933	=>	1548,
		45934	=>	1547,
		45935	=>	1546,
		45936	=>	1545,
		45937	=>	1544,
		45938	=>	1543,
		45939	=>	1542,
		45940	=>	1541,
		45941	=>	1540,
		45942	=>	1540,
		45943	=>	1539,
		45944	=>	1538,
		45945	=>	1537,
		45946	=>	1536,
		45947	=>	1535,
		45948	=>	1534,
		45949	=>	1533,
		45950	=>	1532,
		45951	=>	1531,
		45952	=>	1530,
		45953	=>	1529,
		45954	=>	1528,
		45955	=>	1527,
		45956	=>	1526,
		45957	=>	1525,
		45958	=>	1524,
		45959	=>	1523,
		45960	=>	1522,
		45961	=>	1522,
		45962	=>	1521,
		45963	=>	1520,
		45964	=>	1519,
		45965	=>	1518,
		45966	=>	1517,
		45967	=>	1516,
		45968	=>	1515,
		45969	=>	1514,
		45970	=>	1513,
		45971	=>	1512,
		45972	=>	1511,
		45973	=>	1510,
		45974	=>	1509,
		45975	=>	1508,
		45976	=>	1507,
		45977	=>	1506,
		45978	=>	1505,
		45979	=>	1505,
		45980	=>	1504,
		45981	=>	1503,
		45982	=>	1502,
		45983	=>	1501,
		45984	=>	1500,
		45985	=>	1499,
		45986	=>	1498,
		45987	=>	1497,
		45988	=>	1496,
		45989	=>	1495,
		45990	=>	1494,
		45991	=>	1493,
		45992	=>	1492,
		45993	=>	1491,
		45994	=>	1490,
		45995	=>	1490,
		45996	=>	1489,
		45997	=>	1488,
		45998	=>	1487,
		45999	=>	1486,
		46000	=>	1485,
		46001	=>	1484,
		46002	=>	1483,
		46003	=>	1482,
		46004	=>	1481,
		46005	=>	1480,
		46006	=>	1479,
		46007	=>	1478,
		46008	=>	1477,
		46009	=>	1476,
		46010	=>	1475,
		46011	=>	1475,
		46012	=>	1474,
		46013	=>	1473,
		46014	=>	1472,
		46015	=>	1471,
		46016	=>	1470,
		46017	=>	1469,
		46018	=>	1468,
		46019	=>	1467,
		46020	=>	1466,
		46021	=>	1465,
		46022	=>	1464,
		46023	=>	1463,
		46024	=>	1462,
		46025	=>	1462,
		46026	=>	1461,
		46027	=>	1460,
		46028	=>	1459,
		46029	=>	1458,
		46030	=>	1457,
		46031	=>	1456,
		46032	=>	1455,
		46033	=>	1454,
		46034	=>	1453,
		46035	=>	1452,
		46036	=>	1451,
		46037	=>	1450,
		46038	=>	1450,
		46039	=>	1449,
		46040	=>	1448,
		46041	=>	1447,
		46042	=>	1446,
		46043	=>	1445,
		46044	=>	1444,
		46045	=>	1443,
		46046	=>	1442,
		46047	=>	1441,
		46048	=>	1440,
		46049	=>	1439,
		46050	=>	1438,
		46051	=>	1438,
		46052	=>	1437,
		46053	=>	1436,
		46054	=>	1435,
		46055	=>	1434,
		46056	=>	1433,
		46057	=>	1432,
		46058	=>	1431,
		46059	=>	1430,
		46060	=>	1429,
		46061	=>	1428,
		46062	=>	1427,
		46063	=>	1427,
		46064	=>	1426,
		46065	=>	1425,
		46066	=>	1424,
		46067	=>	1423,
		46068	=>	1422,
		46069	=>	1421,
		46070	=>	1420,
		46071	=>	1419,
		46072	=>	1418,
		46073	=>	1417,
		46074	=>	1416,
		46075	=>	1416,
		46076	=>	1415,
		46077	=>	1414,
		46078	=>	1413,
		46079	=>	1412,
		46080	=>	1411,
		46081	=>	1410,
		46082	=>	1409,
		46083	=>	1408,
		46084	=>	1407,
		46085	=>	1406,
		46086	=>	1405,
		46087	=>	1405,
		46088	=>	1404,
		46089	=>	1403,
		46090	=>	1402,
		46091	=>	1401,
		46092	=>	1400,
		46093	=>	1399,
		46094	=>	1398,
		46095	=>	1397,
		46096	=>	1396,
		46097	=>	1395,
		46098	=>	1395,
		46099	=>	1394,
		46100	=>	1393,
		46101	=>	1392,
		46102	=>	1391,
		46103	=>	1390,
		46104	=>	1389,
		46105	=>	1388,
		46106	=>	1387,
		46107	=>	1386,
		46108	=>	1386,
		46109	=>	1385,
		46110	=>	1384,
		46111	=>	1383,
		46112	=>	1382,
		46113	=>	1381,
		46114	=>	1380,
		46115	=>	1379,
		46116	=>	1378,
		46117	=>	1377,
		46118	=>	1377,
		46119	=>	1376,
		46120	=>	1375,
		46121	=>	1374,
		46122	=>	1373,
		46123	=>	1372,
		46124	=>	1371,
		46125	=>	1370,
		46126	=>	1369,
		46127	=>	1368,
		46128	=>	1368,
		46129	=>	1367,
		46130	=>	1366,
		46131	=>	1365,
		46132	=>	1364,
		46133	=>	1363,
		46134	=>	1362,
		46135	=>	1361,
		46136	=>	1360,
		46137	=>	1359,
		46138	=>	1359,
		46139	=>	1358,
		46140	=>	1357,
		46141	=>	1356,
		46142	=>	1355,
		46143	=>	1354,
		46144	=>	1353,
		46145	=>	1352,
		46146	=>	1351,
		46147	=>	1351,
		46148	=>	1350,
		46149	=>	1349,
		46150	=>	1348,
		46151	=>	1347,
		46152	=>	1346,
		46153	=>	1345,
		46154	=>	1344,
		46155	=>	1343,
		46156	=>	1342,
		46157	=>	1342,
		46158	=>	1341,
		46159	=>	1340,
		46160	=>	1339,
		46161	=>	1338,
		46162	=>	1337,
		46163	=>	1336,
		46164	=>	1335,
		46165	=>	1334,
		46166	=>	1334,
		46167	=>	1333,
		46168	=>	1332,
		46169	=>	1331,
		46170	=>	1330,
		46171	=>	1329,
		46172	=>	1328,
		46173	=>	1327,
		46174	=>	1327,
		46175	=>	1326,
		46176	=>	1325,
		46177	=>	1324,
		46178	=>	1323,
		46179	=>	1322,
		46180	=>	1321,
		46181	=>	1320,
		46182	=>	1319,
		46183	=>	1319,
		46184	=>	1318,
		46185	=>	1317,
		46186	=>	1316,
		46187	=>	1315,
		46188	=>	1314,
		46189	=>	1313,
		46190	=>	1312,
		46191	=>	1312,
		46192	=>	1311,
		46193	=>	1310,
		46194	=>	1309,
		46195	=>	1308,
		46196	=>	1307,
		46197	=>	1306,
		46198	=>	1305,
		46199	=>	1304,
		46200	=>	1304,
		46201	=>	1303,
		46202	=>	1302,
		46203	=>	1301,
		46204	=>	1300,
		46205	=>	1299,
		46206	=>	1298,
		46207	=>	1297,
		46208	=>	1297,
		46209	=>	1296,
		46210	=>	1295,
		46211	=>	1294,
		46212	=>	1293,
		46213	=>	1292,
		46214	=>	1291,
		46215	=>	1290,
		46216	=>	1290,
		46217	=>	1289,
		46218	=>	1288,
		46219	=>	1287,
		46220	=>	1286,
		46221	=>	1285,
		46222	=>	1284,
		46223	=>	1284,
		46224	=>	1283,
		46225	=>	1282,
		46226	=>	1281,
		46227	=>	1280,
		46228	=>	1279,
		46229	=>	1278,
		46230	=>	1277,
		46231	=>	1277,
		46232	=>	1276,
		46233	=>	1275,
		46234	=>	1274,
		46235	=>	1273,
		46236	=>	1272,
		46237	=>	1271,
		46238	=>	1270,
		46239	=>	1270,
		46240	=>	1269,
		46241	=>	1268,
		46242	=>	1267,
		46243	=>	1266,
		46244	=>	1265,
		46245	=>	1264,
		46246	=>	1264,
		46247	=>	1263,
		46248	=>	1262,
		46249	=>	1261,
		46250	=>	1260,
		46251	=>	1259,
		46252	=>	1258,
		46253	=>	1258,
		46254	=>	1257,
		46255	=>	1256,
		46256	=>	1255,
		46257	=>	1254,
		46258	=>	1253,
		46259	=>	1252,
		46260	=>	1251,
		46261	=>	1251,
		46262	=>	1250,
		46263	=>	1249,
		46264	=>	1248,
		46265	=>	1247,
		46266	=>	1246,
		46267	=>	1245,
		46268	=>	1245,
		46269	=>	1244,
		46270	=>	1243,
		46271	=>	1242,
		46272	=>	1241,
		46273	=>	1240,
		46274	=>	1239,
		46275	=>	1239,
		46276	=>	1238,
		46277	=>	1237,
		46278	=>	1236,
		46279	=>	1235,
		46280	=>	1234,
		46281	=>	1233,
		46282	=>	1233,
		46283	=>	1232,
		46284	=>	1231,
		46285	=>	1230,
		46286	=>	1229,
		46287	=>	1228,
		46288	=>	1228,
		46289	=>	1227,
		46290	=>	1226,
		46291	=>	1225,
		46292	=>	1224,
		46293	=>	1223,
		46294	=>	1222,
		46295	=>	1222,
		46296	=>	1221,
		46297	=>	1220,
		46298	=>	1219,
		46299	=>	1218,
		46300	=>	1217,
		46301	=>	1216,
		46302	=>	1216,
		46303	=>	1215,
		46304	=>	1214,
		46305	=>	1213,
		46306	=>	1212,
		46307	=>	1211,
		46308	=>	1211,
		46309	=>	1210,
		46310	=>	1209,
		46311	=>	1208,
		46312	=>	1207,
		46313	=>	1206,
		46314	=>	1205,
		46315	=>	1205,
		46316	=>	1204,
		46317	=>	1203,
		46318	=>	1202,
		46319	=>	1201,
		46320	=>	1200,
		46321	=>	1200,
		46322	=>	1199,
		46323	=>	1198,
		46324	=>	1197,
		46325	=>	1196,
		46326	=>	1195,
		46327	=>	1195,
		46328	=>	1194,
		46329	=>	1193,
		46330	=>	1192,
		46331	=>	1191,
		46332	=>	1190,
		46333	=>	1189,
		46334	=>	1189,
		46335	=>	1188,
		46336	=>	1187,
		46337	=>	1186,
		46338	=>	1185,
		46339	=>	1184,
		46340	=>	1184,
		46341	=>	1183,
		46342	=>	1182,
		46343	=>	1181,
		46344	=>	1180,
		46345	=>	1179,
		46346	=>	1179,
		46347	=>	1178,
		46348	=>	1177,
		46349	=>	1176,
		46350	=>	1175,
		46351	=>	1174,
		46352	=>	1174,
		46353	=>	1173,
		46354	=>	1172,
		46355	=>	1171,
		46356	=>	1170,
		46357	=>	1169,
		46358	=>	1169,
		46359	=>	1168,
		46360	=>	1167,
		46361	=>	1166,
		46362	=>	1165,
		46363	=>	1164,
		46364	=>	1164,
		46365	=>	1163,
		46366	=>	1162,
		46367	=>	1161,
		46368	=>	1160,
		46369	=>	1159,
		46370	=>	1159,
		46371	=>	1158,
		46372	=>	1157,
		46373	=>	1156,
		46374	=>	1155,
		46375	=>	1155,
		46376	=>	1154,
		46377	=>	1153,
		46378	=>	1152,
		46379	=>	1151,
		46380	=>	1150,
		46381	=>	1150,
		46382	=>	1149,
		46383	=>	1148,
		46384	=>	1147,
		46385	=>	1146,
		46386	=>	1145,
		46387	=>	1145,
		46388	=>	1144,
		46389	=>	1143,
		46390	=>	1142,
		46391	=>	1141,
		46392	=>	1141,
		46393	=>	1140,
		46394	=>	1139,
		46395	=>	1138,
		46396	=>	1137,
		46397	=>	1136,
		46398	=>	1136,
		46399	=>	1135,
		46400	=>	1134,
		46401	=>	1133,
		46402	=>	1132,
		46403	=>	1131,
		46404	=>	1131,
		46405	=>	1130,
		46406	=>	1129,
		46407	=>	1128,
		46408	=>	1127,
		46409	=>	1127,
		46410	=>	1126,
		46411	=>	1125,
		46412	=>	1124,
		46413	=>	1123,
		46414	=>	1122,
		46415	=>	1122,
		46416	=>	1121,
		46417	=>	1120,
		46418	=>	1119,
		46419	=>	1118,
		46420	=>	1118,
		46421	=>	1117,
		46422	=>	1116,
		46423	=>	1115,
		46424	=>	1114,
		46425	=>	1114,
		46426	=>	1113,
		46427	=>	1112,
		46428	=>	1111,
		46429	=>	1110,
		46430	=>	1109,
		46431	=>	1109,
		46432	=>	1108,
		46433	=>	1107,
		46434	=>	1106,
		46435	=>	1105,
		46436	=>	1105,
		46437	=>	1104,
		46438	=>	1103,
		46439	=>	1102,
		46440	=>	1101,
		46441	=>	1101,
		46442	=>	1100,
		46443	=>	1099,
		46444	=>	1098,
		46445	=>	1097,
		46446	=>	1097,
		46447	=>	1096,
		46448	=>	1095,
		46449	=>	1094,
		46450	=>	1093,
		46451	=>	1093,
		46452	=>	1092,
		46453	=>	1091,
		46454	=>	1090,
		46455	=>	1089,
		46456	=>	1089,
		46457	=>	1088,
		46458	=>	1087,
		46459	=>	1086,
		46460	=>	1085,
		46461	=>	1085,
		46462	=>	1084,
		46463	=>	1083,
		46464	=>	1082,
		46465	=>	1081,
		46466	=>	1080,
		46467	=>	1080,
		46468	=>	1079,
		46469	=>	1078,
		46470	=>	1077,
		46471	=>	1077,
		46472	=>	1076,
		46473	=>	1075,
		46474	=>	1074,
		46475	=>	1073,
		46476	=>	1073,
		46477	=>	1072,
		46478	=>	1071,
		46479	=>	1070,
		46480	=>	1069,
		46481	=>	1069,
		46482	=>	1068,
		46483	=>	1067,
		46484	=>	1066,
		46485	=>	1065,
		46486	=>	1065,
		46487	=>	1064,
		46488	=>	1063,
		46489	=>	1062,
		46490	=>	1061,
		46491	=>	1061,
		46492	=>	1060,
		46493	=>	1059,
		46494	=>	1058,
		46495	=>	1057,
		46496	=>	1057,
		46497	=>	1056,
		46498	=>	1055,
		46499	=>	1054,
		46500	=>	1053,
		46501	=>	1053,
		46502	=>	1052,
		46503	=>	1051,
		46504	=>	1050,
		46505	=>	1050,
		46506	=>	1049,
		46507	=>	1048,
		46508	=>	1047,
		46509	=>	1046,
		46510	=>	1046,
		46511	=>	1045,
		46512	=>	1044,
		46513	=>	1043,
		46514	=>	1042,
		46515	=>	1042,
		46516	=>	1041,
		46517	=>	1040,
		46518	=>	1039,
		46519	=>	1039,
		46520	=>	1038,
		46521	=>	1037,
		46522	=>	1036,
		46523	=>	1035,
		46524	=>	1035,
		46525	=>	1034,
		46526	=>	1033,
		46527	=>	1032,
		46528	=>	1031,
		46529	=>	1031,
		46530	=>	1030,
		46531	=>	1029,
		46532	=>	1028,
		46533	=>	1028,
		46534	=>	1027,
		46535	=>	1026,
		46536	=>	1025,
		46537	=>	1024,
		46538	=>	1024,
		46539	=>	1023,
		46540	=>	1022,
		46541	=>	1021,
		46542	=>	1021,
		46543	=>	1020,
		46544	=>	1019,
		46545	=>	1018,
		46546	=>	1017,
		46547	=>	1017,
		46548	=>	1016,
		46549	=>	1015,
		46550	=>	1014,
		46551	=>	1014,
		46552	=>	1013,
		46553	=>	1012,
		46554	=>	1011,
		46555	=>	1010,
		46556	=>	1010,
		46557	=>	1009,
		46558	=>	1008,
		46559	=>	1007,
		46560	=>	1007,
		46561	=>	1006,
		46562	=>	1005,
		46563	=>	1004,
		46564	=>	1003,
		46565	=>	1003,
		46566	=>	1002,
		46567	=>	1001,
		46568	=>	1000,
		46569	=>	1000,
		46570	=>	999,
		46571	=>	998,
		46572	=>	997,
		46573	=>	997,
		46574	=>	996,
		46575	=>	995,
		46576	=>	994,
		46577	=>	993,
		46578	=>	993,
		46579	=>	992,
		46580	=>	991,
		46581	=>	990,
		46582	=>	990,
		46583	=>	989,
		46584	=>	988,
		46585	=>	987,
		46586	=>	987,
		46587	=>	986,
		46588	=>	985,
		46589	=>	984,
		46590	=>	984,
		46591	=>	983,
		46592	=>	982,
		46593	=>	981,
		46594	=>	980,
		46595	=>	980,
		46596	=>	979,
		46597	=>	978,
		46598	=>	977,
		46599	=>	977,
		46600	=>	976,
		46601	=>	975,
		46602	=>	974,
		46603	=>	974,
		46604	=>	973,
		46605	=>	972,
		46606	=>	971,
		46607	=>	971,
		46608	=>	970,
		46609	=>	969,
		46610	=>	968,
		46611	=>	968,
		46612	=>	967,
		46613	=>	966,
		46614	=>	965,
		46615	=>	965,
		46616	=>	964,
		46617	=>	963,
		46618	=>	962,
		46619	=>	961,
		46620	=>	961,
		46621	=>	960,
		46622	=>	959,
		46623	=>	958,
		46624	=>	958,
		46625	=>	957,
		46626	=>	956,
		46627	=>	955,
		46628	=>	955,
		46629	=>	954,
		46630	=>	953,
		46631	=>	952,
		46632	=>	952,
		46633	=>	951,
		46634	=>	950,
		46635	=>	949,
		46636	=>	949,
		46637	=>	948,
		46638	=>	947,
		46639	=>	946,
		46640	=>	946,
		46641	=>	945,
		46642	=>	944,
		46643	=>	943,
		46644	=>	943,
		46645	=>	942,
		46646	=>	941,
		46647	=>	940,
		46648	=>	940,
		46649	=>	939,
		46650	=>	938,
		46651	=>	937,
		46652	=>	937,
		46653	=>	936,
		46654	=>	935,
		46655	=>	934,
		46656	=>	934,
		46657	=>	933,
		46658	=>	932,
		46659	=>	932,
		46660	=>	931,
		46661	=>	930,
		46662	=>	929,
		46663	=>	929,
		46664	=>	928,
		46665	=>	927,
		46666	=>	926,
		46667	=>	926,
		46668	=>	925,
		46669	=>	924,
		46670	=>	923,
		46671	=>	923,
		46672	=>	922,
		46673	=>	921,
		46674	=>	920,
		46675	=>	920,
		46676	=>	919,
		46677	=>	918,
		46678	=>	917,
		46679	=>	917,
		46680	=>	916,
		46681	=>	915,
		46682	=>	914,
		46683	=>	914,
		46684	=>	913,
		46685	=>	912,
		46686	=>	912,
		46687	=>	911,
		46688	=>	910,
		46689	=>	909,
		46690	=>	909,
		46691	=>	908,
		46692	=>	907,
		46693	=>	906,
		46694	=>	906,
		46695	=>	905,
		46696	=>	904,
		46697	=>	903,
		46698	=>	903,
		46699	=>	902,
		46700	=>	901,
		46701	=>	901,
		46702	=>	900,
		46703	=>	899,
		46704	=>	898,
		46705	=>	898,
		46706	=>	897,
		46707	=>	896,
		46708	=>	895,
		46709	=>	895,
		46710	=>	894,
		46711	=>	893,
		46712	=>	893,
		46713	=>	892,
		46714	=>	891,
		46715	=>	890,
		46716	=>	890,
		46717	=>	889,
		46718	=>	888,
		46719	=>	887,
		46720	=>	887,
		46721	=>	886,
		46722	=>	885,
		46723	=>	885,
		46724	=>	884,
		46725	=>	883,
		46726	=>	882,
		46727	=>	882,
		46728	=>	881,
		46729	=>	880,
		46730	=>	879,
		46731	=>	879,
		46732	=>	878,
		46733	=>	877,
		46734	=>	877,
		46735	=>	876,
		46736	=>	875,
		46737	=>	874,
		46738	=>	874,
		46739	=>	873,
		46740	=>	872,
		46741	=>	872,
		46742	=>	871,
		46743	=>	870,
		46744	=>	869,
		46745	=>	869,
		46746	=>	868,
		46747	=>	867,
		46748	=>	866,
		46749	=>	866,
		46750	=>	865,
		46751	=>	864,
		46752	=>	864,
		46753	=>	863,
		46754	=>	862,
		46755	=>	861,
		46756	=>	861,
		46757	=>	860,
		46758	=>	859,
		46759	=>	859,
		46760	=>	858,
		46761	=>	857,
		46762	=>	856,
		46763	=>	856,
		46764	=>	855,
		46765	=>	854,
		46766	=>	854,
		46767	=>	853,
		46768	=>	852,
		46769	=>	851,
		46770	=>	851,
		46771	=>	850,
		46772	=>	849,
		46773	=>	849,
		46774	=>	848,
		46775	=>	847,
		46776	=>	847,
		46777	=>	846,
		46778	=>	845,
		46779	=>	844,
		46780	=>	844,
		46781	=>	843,
		46782	=>	842,
		46783	=>	842,
		46784	=>	841,
		46785	=>	840,
		46786	=>	839,
		46787	=>	839,
		46788	=>	838,
		46789	=>	837,
		46790	=>	837,
		46791	=>	836,
		46792	=>	835,
		46793	=>	834,
		46794	=>	834,
		46795	=>	833,
		46796	=>	832,
		46797	=>	832,
		46798	=>	831,
		46799	=>	830,
		46800	=>	830,
		46801	=>	829,
		46802	=>	828,
		46803	=>	827,
		46804	=>	827,
		46805	=>	826,
		46806	=>	825,
		46807	=>	825,
		46808	=>	824,
		46809	=>	823,
		46810	=>	823,
		46811	=>	822,
		46812	=>	821,
		46813	=>	820,
		46814	=>	820,
		46815	=>	819,
		46816	=>	818,
		46817	=>	818,
		46818	=>	817,
		46819	=>	816,
		46820	=>	816,
		46821	=>	815,
		46822	=>	814,
		46823	=>	813,
		46824	=>	813,
		46825	=>	812,
		46826	=>	811,
		46827	=>	811,
		46828	=>	810,
		46829	=>	809,
		46830	=>	809,
		46831	=>	808,
		46832	=>	807,
		46833	=>	807,
		46834	=>	806,
		46835	=>	805,
		46836	=>	804,
		46837	=>	804,
		46838	=>	803,
		46839	=>	802,
		46840	=>	802,
		46841	=>	801,
		46842	=>	800,
		46843	=>	800,
		46844	=>	799,
		46845	=>	798,
		46846	=>	798,
		46847	=>	797,
		46848	=>	796,
		46849	=>	795,
		46850	=>	795,
		46851	=>	794,
		46852	=>	793,
		46853	=>	793,
		46854	=>	792,
		46855	=>	791,
		46856	=>	791,
		46857	=>	790,
		46858	=>	789,
		46859	=>	789,
		46860	=>	788,
		46861	=>	787,
		46862	=>	787,
		46863	=>	786,
		46864	=>	785,
		46865	=>	785,
		46866	=>	784,
		46867	=>	783,
		46868	=>	782,
		46869	=>	782,
		46870	=>	781,
		46871	=>	780,
		46872	=>	780,
		46873	=>	779,
		46874	=>	778,
		46875	=>	778,
		46876	=>	777,
		46877	=>	776,
		46878	=>	776,
		46879	=>	775,
		46880	=>	774,
		46881	=>	774,
		46882	=>	773,
		46883	=>	772,
		46884	=>	772,
		46885	=>	771,
		46886	=>	770,
		46887	=>	770,
		46888	=>	769,
		46889	=>	768,
		46890	=>	768,
		46891	=>	767,
		46892	=>	766,
		46893	=>	766,
		46894	=>	765,
		46895	=>	764,
		46896	=>	763,
		46897	=>	763,
		46898	=>	762,
		46899	=>	761,
		46900	=>	761,
		46901	=>	760,
		46902	=>	759,
		46903	=>	759,
		46904	=>	758,
		46905	=>	757,
		46906	=>	757,
		46907	=>	756,
		46908	=>	755,
		46909	=>	755,
		46910	=>	754,
		46911	=>	753,
		46912	=>	753,
		46913	=>	752,
		46914	=>	751,
		46915	=>	751,
		46916	=>	750,
		46917	=>	749,
		46918	=>	749,
		46919	=>	748,
		46920	=>	747,
		46921	=>	747,
		46922	=>	746,
		46923	=>	745,
		46924	=>	745,
		46925	=>	744,
		46926	=>	743,
		46927	=>	743,
		46928	=>	742,
		46929	=>	741,
		46930	=>	741,
		46931	=>	740,
		46932	=>	739,
		46933	=>	739,
		46934	=>	738,
		46935	=>	737,
		46936	=>	737,
		46937	=>	736,
		46938	=>	735,
		46939	=>	735,
		46940	=>	734,
		46941	=>	733,
		46942	=>	733,
		46943	=>	732,
		46944	=>	731,
		46945	=>	731,
		46946	=>	730,
		46947	=>	729,
		46948	=>	729,
		46949	=>	728,
		46950	=>	728,
		46951	=>	727,
		46952	=>	726,
		46953	=>	726,
		46954	=>	725,
		46955	=>	724,
		46956	=>	724,
		46957	=>	723,
		46958	=>	722,
		46959	=>	722,
		46960	=>	721,
		46961	=>	720,
		46962	=>	720,
		46963	=>	719,
		46964	=>	718,
		46965	=>	718,
		46966	=>	717,
		46967	=>	716,
		46968	=>	716,
		46969	=>	715,
		46970	=>	714,
		46971	=>	714,
		46972	=>	713,
		46973	=>	712,
		46974	=>	712,
		46975	=>	711,
		46976	=>	710,
		46977	=>	710,
		46978	=>	709,
		46979	=>	709,
		46980	=>	708,
		46981	=>	707,
		46982	=>	707,
		46983	=>	706,
		46984	=>	705,
		46985	=>	705,
		46986	=>	704,
		46987	=>	703,
		46988	=>	703,
		46989	=>	702,
		46990	=>	701,
		46991	=>	701,
		46992	=>	700,
		46993	=>	699,
		46994	=>	699,
		46995	=>	698,
		46996	=>	698,
		46997	=>	697,
		46998	=>	696,
		46999	=>	696,
		47000	=>	695,
		47001	=>	694,
		47002	=>	694,
		47003	=>	693,
		47004	=>	692,
		47005	=>	692,
		47006	=>	691,
		47007	=>	690,
		47008	=>	690,
		47009	=>	689,
		47010	=>	689,
		47011	=>	688,
		47012	=>	687,
		47013	=>	687,
		47014	=>	686,
		47015	=>	685,
		47016	=>	685,
		47017	=>	684,
		47018	=>	683,
		47019	=>	683,
		47020	=>	682,
		47021	=>	682,
		47022	=>	681,
		47023	=>	680,
		47024	=>	680,
		47025	=>	679,
		47026	=>	678,
		47027	=>	678,
		47028	=>	677,
		47029	=>	676,
		47030	=>	676,
		47031	=>	675,
		47032	=>	675,
		47033	=>	674,
		47034	=>	673,
		47035	=>	673,
		47036	=>	672,
		47037	=>	671,
		47038	=>	671,
		47039	=>	670,
		47040	=>	669,
		47041	=>	669,
		47042	=>	668,
		47043	=>	668,
		47044	=>	667,
		47045	=>	666,
		47046	=>	666,
		47047	=>	665,
		47048	=>	664,
		47049	=>	664,
		47050	=>	663,
		47051	=>	663,
		47052	=>	662,
		47053	=>	661,
		47054	=>	661,
		47055	=>	660,
		47056	=>	659,
		47057	=>	659,
		47058	=>	658,
		47059	=>	657,
		47060	=>	657,
		47061	=>	656,
		47062	=>	656,
		47063	=>	655,
		47064	=>	654,
		47065	=>	654,
		47066	=>	653,
		47067	=>	652,
		47068	=>	652,
		47069	=>	651,
		47070	=>	651,
		47071	=>	650,
		47072	=>	649,
		47073	=>	649,
		47074	=>	648,
		47075	=>	648,
		47076	=>	647,
		47077	=>	646,
		47078	=>	646,
		47079	=>	645,
		47080	=>	644,
		47081	=>	644,
		47082	=>	643,
		47083	=>	643,
		47084	=>	642,
		47085	=>	641,
		47086	=>	641,
		47087	=>	640,
		47088	=>	639,
		47089	=>	639,
		47090	=>	638,
		47091	=>	638,
		47092	=>	637,
		47093	=>	636,
		47094	=>	636,
		47095	=>	635,
		47096	=>	635,
		47097	=>	634,
		47098	=>	633,
		47099	=>	633,
		47100	=>	632,
		47101	=>	631,
		47102	=>	631,
		47103	=>	630,
		47104	=>	630,
		47105	=>	629,
		47106	=>	628,
		47107	=>	628,
		47108	=>	627,
		47109	=>	627,
		47110	=>	626,
		47111	=>	625,
		47112	=>	625,
		47113	=>	624,
		47114	=>	624,
		47115	=>	623,
		47116	=>	622,
		47117	=>	622,
		47118	=>	621,
		47119	=>	620,
		47120	=>	620,
		47121	=>	619,
		47122	=>	619,
		47123	=>	618,
		47124	=>	617,
		47125	=>	617,
		47126	=>	616,
		47127	=>	616,
		47128	=>	615,
		47129	=>	614,
		47130	=>	614,
		47131	=>	613,
		47132	=>	613,
		47133	=>	612,
		47134	=>	611,
		47135	=>	611,
		47136	=>	610,
		47137	=>	610,
		47138	=>	609,
		47139	=>	608,
		47140	=>	608,
		47141	=>	607,
		47142	=>	607,
		47143	=>	606,
		47144	=>	605,
		47145	=>	605,
		47146	=>	604,
		47147	=>	604,
		47148	=>	603,
		47149	=>	602,
		47150	=>	602,
		47151	=>	601,
		47152	=>	601,
		47153	=>	600,
		47154	=>	599,
		47155	=>	599,
		47156	=>	598,
		47157	=>	598,
		47158	=>	597,
		47159	=>	596,
		47160	=>	596,
		47161	=>	595,
		47162	=>	595,
		47163	=>	594,
		47164	=>	593,
		47165	=>	593,
		47166	=>	592,
		47167	=>	592,
		47168	=>	591,
		47169	=>	590,
		47170	=>	590,
		47171	=>	589,
		47172	=>	589,
		47173	=>	588,
		47174	=>	587,
		47175	=>	587,
		47176	=>	586,
		47177	=>	586,
		47178	=>	585,
		47179	=>	584,
		47180	=>	584,
		47181	=>	583,
		47182	=>	583,
		47183	=>	582,
		47184	=>	582,
		47185	=>	581,
		47186	=>	580,
		47187	=>	580,
		47188	=>	579,
		47189	=>	579,
		47190	=>	578,
		47191	=>	577,
		47192	=>	577,
		47193	=>	576,
		47194	=>	576,
		47195	=>	575,
		47196	=>	574,
		47197	=>	574,
		47198	=>	573,
		47199	=>	573,
		47200	=>	572,
		47201	=>	572,
		47202	=>	571,
		47203	=>	570,
		47204	=>	570,
		47205	=>	569,
		47206	=>	569,
		47207	=>	568,
		47208	=>	567,
		47209	=>	567,
		47210	=>	566,
		47211	=>	566,
		47212	=>	565,
		47213	=>	565,
		47214	=>	564,
		47215	=>	563,
		47216	=>	563,
		47217	=>	562,
		47218	=>	562,
		47219	=>	561,
		47220	=>	561,
		47221	=>	560,
		47222	=>	559,
		47223	=>	559,
		47224	=>	558,
		47225	=>	558,
		47226	=>	557,
		47227	=>	556,
		47228	=>	556,
		47229	=>	555,
		47230	=>	555,
		47231	=>	554,
		47232	=>	554,
		47233	=>	553,
		47234	=>	552,
		47235	=>	552,
		47236	=>	551,
		47237	=>	551,
		47238	=>	550,
		47239	=>	550,
		47240	=>	549,
		47241	=>	548,
		47242	=>	548,
		47243	=>	547,
		47244	=>	547,
		47245	=>	546,
		47246	=>	546,
		47247	=>	545,
		47248	=>	544,
		47249	=>	544,
		47250	=>	543,
		47251	=>	543,
		47252	=>	542,
		47253	=>	542,
		47254	=>	541,
		47255	=>	540,
		47256	=>	540,
		47257	=>	539,
		47258	=>	539,
		47259	=>	538,
		47260	=>	538,
		47261	=>	537,
		47262	=>	536,
		47263	=>	536,
		47264	=>	535,
		47265	=>	535,
		47266	=>	534,
		47267	=>	534,
		47268	=>	533,
		47269	=>	533,
		47270	=>	532,
		47271	=>	531,
		47272	=>	531,
		47273	=>	530,
		47274	=>	530,
		47275	=>	529,
		47276	=>	529,
		47277	=>	528,
		47278	=>	527,
		47279	=>	527,
		47280	=>	526,
		47281	=>	526,
		47282	=>	525,
		47283	=>	525,
		47284	=>	524,
		47285	=>	524,
		47286	=>	523,
		47287	=>	522,
		47288	=>	522,
		47289	=>	521,
		47290	=>	521,
		47291	=>	520,
		47292	=>	520,
		47293	=>	519,
		47294	=>	519,
		47295	=>	518,
		47296	=>	517,
		47297	=>	517,
		47298	=>	516,
		47299	=>	516,
		47300	=>	515,
		47301	=>	515,
		47302	=>	514,
		47303	=>	514,
		47304	=>	513,
		47305	=>	512,
		47306	=>	512,
		47307	=>	511,
		47308	=>	511,
		47309	=>	510,
		47310	=>	510,
		47311	=>	509,
		47312	=>	509,
		47313	=>	508,
		47314	=>	507,
		47315	=>	507,
		47316	=>	506,
		47317	=>	506,
		47318	=>	505,
		47319	=>	505,
		47320	=>	504,
		47321	=>	504,
		47322	=>	503,
		47323	=>	502,
		47324	=>	502,
		47325	=>	501,
		47326	=>	501,
		47327	=>	500,
		47328	=>	500,
		47329	=>	499,
		47330	=>	499,
		47331	=>	498,
		47332	=>	498,
		47333	=>	497,
		47334	=>	496,
		47335	=>	496,
		47336	=>	495,
		47337	=>	495,
		47338	=>	494,
		47339	=>	494,
		47340	=>	493,
		47341	=>	493,
		47342	=>	492,
		47343	=>	492,
		47344	=>	491,
		47345	=>	491,
		47346	=>	490,
		47347	=>	489,
		47348	=>	489,
		47349	=>	488,
		47350	=>	488,
		47351	=>	487,
		47352	=>	487,
		47353	=>	486,
		47354	=>	486,
		47355	=>	485,
		47356	=>	485,
		47357	=>	484,
		47358	=>	483,
		47359	=>	483,
		47360	=>	482,
		47361	=>	482,
		47362	=>	481,
		47363	=>	481,
		47364	=>	480,
		47365	=>	480,
		47366	=>	479,
		47367	=>	479,
		47368	=>	478,
		47369	=>	478,
		47370	=>	477,
		47371	=>	477,
		47372	=>	476,
		47373	=>	475,
		47374	=>	475,
		47375	=>	474,
		47376	=>	474,
		47377	=>	473,
		47378	=>	473,
		47379	=>	472,
		47380	=>	472,
		47381	=>	471,
		47382	=>	471,
		47383	=>	470,
		47384	=>	470,
		47385	=>	469,
		47386	=>	469,
		47387	=>	468,
		47388	=>	467,
		47389	=>	467,
		47390	=>	466,
		47391	=>	466,
		47392	=>	465,
		47393	=>	465,
		47394	=>	464,
		47395	=>	464,
		47396	=>	463,
		47397	=>	463,
		47398	=>	462,
		47399	=>	462,
		47400	=>	461,
		47401	=>	461,
		47402	=>	460,
		47403	=>	460,
		47404	=>	459,
		47405	=>	459,
		47406	=>	458,
		47407	=>	457,
		47408	=>	457,
		47409	=>	456,
		47410	=>	456,
		47411	=>	455,
		47412	=>	455,
		47413	=>	454,
		47414	=>	454,
		47415	=>	453,
		47416	=>	453,
		47417	=>	452,
		47418	=>	452,
		47419	=>	451,
		47420	=>	451,
		47421	=>	450,
		47422	=>	450,
		47423	=>	449,
		47424	=>	449,
		47425	=>	448,
		47426	=>	448,
		47427	=>	447,
		47428	=>	447,
		47429	=>	446,
		47430	=>	446,
		47431	=>	445,
		47432	=>	445,
		47433	=>	444,
		47434	=>	443,
		47435	=>	443,
		47436	=>	442,
		47437	=>	442,
		47438	=>	441,
		47439	=>	441,
		47440	=>	440,
		47441	=>	440,
		47442	=>	439,
		47443	=>	439,
		47444	=>	438,
		47445	=>	438,
		47446	=>	437,
		47447	=>	437,
		47448	=>	436,
		47449	=>	436,
		47450	=>	435,
		47451	=>	435,
		47452	=>	434,
		47453	=>	434,
		47454	=>	433,
		47455	=>	433,
		47456	=>	432,
		47457	=>	432,
		47458	=>	431,
		47459	=>	431,
		47460	=>	430,
		47461	=>	430,
		47462	=>	429,
		47463	=>	429,
		47464	=>	428,
		47465	=>	428,
		47466	=>	427,
		47467	=>	427,
		47468	=>	426,
		47469	=>	426,
		47470	=>	425,
		47471	=>	425,
		47472	=>	424,
		47473	=>	424,
		47474	=>	423,
		47475	=>	423,
		47476	=>	422,
		47477	=>	422,
		47478	=>	421,
		47479	=>	421,
		47480	=>	420,
		47481	=>	420,
		47482	=>	419,
		47483	=>	419,
		47484	=>	418,
		47485	=>	418,
		47486	=>	417,
		47487	=>	417,
		47488	=>	416,
		47489	=>	416,
		47490	=>	415,
		47491	=>	415,
		47492	=>	414,
		47493	=>	414,
		47494	=>	413,
		47495	=>	413,
		47496	=>	412,
		47497	=>	412,
		47498	=>	411,
		47499	=>	411,
		47500	=>	410,
		47501	=>	410,
		47502	=>	409,
		47503	=>	409,
		47504	=>	408,
		47505	=>	408,
		47506	=>	407,
		47507	=>	407,
		47508	=>	406,
		47509	=>	406,
		47510	=>	405,
		47511	=>	405,
		47512	=>	404,
		47513	=>	404,
		47514	=>	403,
		47515	=>	403,
		47516	=>	402,
		47517	=>	402,
		47518	=>	401,
		47519	=>	401,
		47520	=>	400,
		47521	=>	400,
		47522	=>	399,
		47523	=>	399,
		47524	=>	398,
		47525	=>	398,
		47526	=>	397,
		47527	=>	397,
		47528	=>	396,
		47529	=>	396,
		47530	=>	395,
		47531	=>	395,
		47532	=>	394,
		47533	=>	394,
		47534	=>	393,
		47535	=>	393,
		47536	=>	392,
		47537	=>	392,
		47538	=>	392,
		47539	=>	391,
		47540	=>	391,
		47541	=>	390,
		47542	=>	390,
		47543	=>	389,
		47544	=>	389,
		47545	=>	388,
		47546	=>	388,
		47547	=>	387,
		47548	=>	387,
		47549	=>	386,
		47550	=>	386,
		47551	=>	385,
		47552	=>	385,
		47553	=>	384,
		47554	=>	384,
		47555	=>	383,
		47556	=>	383,
		47557	=>	382,
		47558	=>	382,
		47559	=>	381,
		47560	=>	381,
		47561	=>	380,
		47562	=>	380,
		47563	=>	380,
		47564	=>	379,
		47565	=>	379,
		47566	=>	378,
		47567	=>	378,
		47568	=>	377,
		47569	=>	377,
		47570	=>	376,
		47571	=>	376,
		47572	=>	375,
		47573	=>	375,
		47574	=>	374,
		47575	=>	374,
		47576	=>	373,
		47577	=>	373,
		47578	=>	372,
		47579	=>	372,
		47580	=>	371,
		47581	=>	371,
		47582	=>	371,
		47583	=>	370,
		47584	=>	370,
		47585	=>	369,
		47586	=>	369,
		47587	=>	368,
		47588	=>	368,
		47589	=>	367,
		47590	=>	367,
		47591	=>	366,
		47592	=>	366,
		47593	=>	365,
		47594	=>	365,
		47595	=>	364,
		47596	=>	364,
		47597	=>	363,
		47598	=>	363,
		47599	=>	363,
		47600	=>	362,
		47601	=>	362,
		47602	=>	361,
		47603	=>	361,
		47604	=>	360,
		47605	=>	360,
		47606	=>	359,
		47607	=>	359,
		47608	=>	358,
		47609	=>	358,
		47610	=>	357,
		47611	=>	357,
		47612	=>	357,
		47613	=>	356,
		47614	=>	356,
		47615	=>	355,
		47616	=>	355,
		47617	=>	354,
		47618	=>	354,
		47619	=>	353,
		47620	=>	353,
		47621	=>	352,
		47622	=>	352,
		47623	=>	351,
		47624	=>	351,
		47625	=>	351,
		47626	=>	350,
		47627	=>	350,
		47628	=>	349,
		47629	=>	349,
		47630	=>	348,
		47631	=>	348,
		47632	=>	347,
		47633	=>	347,
		47634	=>	346,
		47635	=>	346,
		47636	=>	345,
		47637	=>	345,
		47638	=>	345,
		47639	=>	344,
		47640	=>	344,
		47641	=>	343,
		47642	=>	343,
		47643	=>	342,
		47644	=>	342,
		47645	=>	341,
		47646	=>	341,
		47647	=>	341,
		47648	=>	340,
		47649	=>	340,
		47650	=>	339,
		47651	=>	339,
		47652	=>	338,
		47653	=>	338,
		47654	=>	337,
		47655	=>	337,
		47656	=>	336,
		47657	=>	336,
		47658	=>	336,
		47659	=>	335,
		47660	=>	335,
		47661	=>	334,
		47662	=>	334,
		47663	=>	333,
		47664	=>	333,
		47665	=>	332,
		47666	=>	332,
		47667	=>	332,
		47668	=>	331,
		47669	=>	331,
		47670	=>	330,
		47671	=>	330,
		47672	=>	329,
		47673	=>	329,
		47674	=>	328,
		47675	=>	328,
		47676	=>	328,
		47677	=>	327,
		47678	=>	327,
		47679	=>	326,
		47680	=>	326,
		47681	=>	325,
		47682	=>	325,
		47683	=>	324,
		47684	=>	324,
		47685	=>	324,
		47686	=>	323,
		47687	=>	323,
		47688	=>	322,
		47689	=>	322,
		47690	=>	321,
		47691	=>	321,
		47692	=>	320,
		47693	=>	320,
		47694	=>	320,
		47695	=>	319,
		47696	=>	319,
		47697	=>	318,
		47698	=>	318,
		47699	=>	317,
		47700	=>	317,
		47701	=>	317,
		47702	=>	316,
		47703	=>	316,
		47704	=>	315,
		47705	=>	315,
		47706	=>	314,
		47707	=>	314,
		47708	=>	314,
		47709	=>	313,
		47710	=>	313,
		47711	=>	312,
		47712	=>	312,
		47713	=>	311,
		47714	=>	311,
		47715	=>	310,
		47716	=>	310,
		47717	=>	310,
		47718	=>	309,
		47719	=>	309,
		47720	=>	308,
		47721	=>	308,
		47722	=>	307,
		47723	=>	307,
		47724	=>	307,
		47725	=>	306,
		47726	=>	306,
		47727	=>	305,
		47728	=>	305,
		47729	=>	304,
		47730	=>	304,
		47731	=>	304,
		47732	=>	303,
		47733	=>	303,
		47734	=>	302,
		47735	=>	302,
		47736	=>	301,
		47737	=>	301,
		47738	=>	301,
		47739	=>	300,
		47740	=>	300,
		47741	=>	299,
		47742	=>	299,
		47743	=>	299,
		47744	=>	298,
		47745	=>	298,
		47746	=>	297,
		47747	=>	297,
		47748	=>	296,
		47749	=>	296,
		47750	=>	296,
		47751	=>	295,
		47752	=>	295,
		47753	=>	294,
		47754	=>	294,
		47755	=>	293,
		47756	=>	293,
		47757	=>	293,
		47758	=>	292,
		47759	=>	292,
		47760	=>	291,
		47761	=>	291,
		47762	=>	291,
		47763	=>	290,
		47764	=>	290,
		47765	=>	289,
		47766	=>	289,
		47767	=>	288,
		47768	=>	288,
		47769	=>	288,
		47770	=>	287,
		47771	=>	287,
		47772	=>	286,
		47773	=>	286,
		47774	=>	286,
		47775	=>	285,
		47776	=>	285,
		47777	=>	284,
		47778	=>	284,
		47779	=>	283,
		47780	=>	283,
		47781	=>	283,
		47782	=>	282,
		47783	=>	282,
		47784	=>	281,
		47785	=>	281,
		47786	=>	281,
		47787	=>	280,
		47788	=>	280,
		47789	=>	279,
		47790	=>	279,
		47791	=>	279,
		47792	=>	278,
		47793	=>	278,
		47794	=>	277,
		47795	=>	277,
		47796	=>	277,
		47797	=>	276,
		47798	=>	276,
		47799	=>	275,
		47800	=>	275,
		47801	=>	274,
		47802	=>	274,
		47803	=>	274,
		47804	=>	273,
		47805	=>	273,
		47806	=>	272,
		47807	=>	272,
		47808	=>	272,
		47809	=>	271,
		47810	=>	271,
		47811	=>	270,
		47812	=>	270,
		47813	=>	270,
		47814	=>	269,
		47815	=>	269,
		47816	=>	268,
		47817	=>	268,
		47818	=>	268,
		47819	=>	267,
		47820	=>	267,
		47821	=>	266,
		47822	=>	266,
		47823	=>	266,
		47824	=>	265,
		47825	=>	265,
		47826	=>	264,
		47827	=>	264,
		47828	=>	264,
		47829	=>	263,
		47830	=>	263,
		47831	=>	262,
		47832	=>	262,
		47833	=>	262,
		47834	=>	261,
		47835	=>	261,
		47836	=>	260,
		47837	=>	260,
		47838	=>	260,
		47839	=>	259,
		47840	=>	259,
		47841	=>	258,
		47842	=>	258,
		47843	=>	258,
		47844	=>	257,
		47845	=>	257,
		47846	=>	257,
		47847	=>	256,
		47848	=>	256,
		47849	=>	255,
		47850	=>	255,
		47851	=>	255,
		47852	=>	254,
		47853	=>	254,
		47854	=>	253,
		47855	=>	253,
		47856	=>	253,
		47857	=>	252,
		47858	=>	252,
		47859	=>	251,
		47860	=>	251,
		47861	=>	251,
		47862	=>	250,
		47863	=>	250,
		47864	=>	250,
		47865	=>	249,
		47866	=>	249,
		47867	=>	248,
		47868	=>	248,
		47869	=>	248,
		47870	=>	247,
		47871	=>	247,
		47872	=>	246,
		47873	=>	246,
		47874	=>	246,
		47875	=>	245,
		47876	=>	245,
		47877	=>	245,
		47878	=>	244,
		47879	=>	244,
		47880	=>	243,
		47881	=>	243,
		47882	=>	243,
		47883	=>	242,
		47884	=>	242,
		47885	=>	241,
		47886	=>	241,
		47887	=>	241,
		47888	=>	240,
		47889	=>	240,
		47890	=>	240,
		47891	=>	239,
		47892	=>	239,
		47893	=>	238,
		47894	=>	238,
		47895	=>	238,
		47896	=>	237,
		47897	=>	237,
		47898	=>	237,
		47899	=>	236,
		47900	=>	236,
		47901	=>	235,
		47902	=>	235,
		47903	=>	235,
		47904	=>	234,
		47905	=>	234,
		47906	=>	234,
		47907	=>	233,
		47908	=>	233,
		47909	=>	232,
		47910	=>	232,
		47911	=>	232,
		47912	=>	231,
		47913	=>	231,
		47914	=>	231,
		47915	=>	230,
		47916	=>	230,
		47917	=>	229,
		47918	=>	229,
		47919	=>	229,
		47920	=>	228,
		47921	=>	228,
		47922	=>	228,
		47923	=>	227,
		47924	=>	227,
		47925	=>	226,
		47926	=>	226,
		47927	=>	226,
		47928	=>	225,
		47929	=>	225,
		47930	=>	225,
		47931	=>	224,
		47932	=>	224,
		47933	=>	224,
		47934	=>	223,
		47935	=>	223,
		47936	=>	222,
		47937	=>	222,
		47938	=>	222,
		47939	=>	221,
		47940	=>	221,
		47941	=>	221,
		47942	=>	220,
		47943	=>	220,
		47944	=>	220,
		47945	=>	219,
		47946	=>	219,
		47947	=>	218,
		47948	=>	218,
		47949	=>	218,
		47950	=>	217,
		47951	=>	217,
		47952	=>	217,
		47953	=>	216,
		47954	=>	216,
		47955	=>	216,
		47956	=>	215,
		47957	=>	215,
		47958	=>	214,
		47959	=>	214,
		47960	=>	214,
		47961	=>	213,
		47962	=>	213,
		47963	=>	213,
		47964	=>	212,
		47965	=>	212,
		47966	=>	212,
		47967	=>	211,
		47968	=>	211,
		47969	=>	211,
		47970	=>	210,
		47971	=>	210,
		47972	=>	209,
		47973	=>	209,
		47974	=>	209,
		47975	=>	208,
		47976	=>	208,
		47977	=>	208,
		47978	=>	207,
		47979	=>	207,
		47980	=>	207,
		47981	=>	206,
		47982	=>	206,
		47983	=>	206,
		47984	=>	205,
		47985	=>	205,
		47986	=>	205,
		47987	=>	204,
		47988	=>	204,
		47989	=>	203,
		47990	=>	203,
		47991	=>	203,
		47992	=>	202,
		47993	=>	202,
		47994	=>	202,
		47995	=>	201,
		47996	=>	201,
		47997	=>	201,
		47998	=>	200,
		47999	=>	200,
		48000	=>	200,
		48001	=>	199,
		48002	=>	199,
		48003	=>	199,
		48004	=>	198,
		48005	=>	198,
		48006	=>	198,
		48007	=>	197,
		48008	=>	197,
		48009	=>	197,
		48010	=>	196,
		48011	=>	196,
		48012	=>	196,
		48013	=>	195,
		48014	=>	195,
		48015	=>	194,
		48016	=>	194,
		48017	=>	194,
		48018	=>	193,
		48019	=>	193,
		48020	=>	193,
		48021	=>	192,
		48022	=>	192,
		48023	=>	192,
		48024	=>	191,
		48025	=>	191,
		48026	=>	191,
		48027	=>	190,
		48028	=>	190,
		48029	=>	190,
		48030	=>	189,
		48031	=>	189,
		48032	=>	189,
		48033	=>	188,
		48034	=>	188,
		48035	=>	188,
		48036	=>	187,
		48037	=>	187,
		48038	=>	187,
		48039	=>	186,
		48040	=>	186,
		48041	=>	186,
		48042	=>	185,
		48043	=>	185,
		48044	=>	185,
		48045	=>	184,
		48046	=>	184,
		48047	=>	184,
		48048	=>	183,
		48049	=>	183,
		48050	=>	183,
		48051	=>	182,
		48052	=>	182,
		48053	=>	182,
		48054	=>	181,
		48055	=>	181,
		48056	=>	181,
		48057	=>	180,
		48058	=>	180,
		48059	=>	180,
		48060	=>	179,
		48061	=>	179,
		48062	=>	179,
		48063	=>	178,
		48064	=>	178,
		48065	=>	178,
		48066	=>	177,
		48067	=>	177,
		48068	=>	177,
		48069	=>	176,
		48070	=>	176,
		48071	=>	176,
		48072	=>	175,
		48073	=>	175,
		48074	=>	175,
		48075	=>	175,
		48076	=>	174,
		48077	=>	174,
		48078	=>	174,
		48079	=>	173,
		48080	=>	173,
		48081	=>	173,
		48082	=>	172,
		48083	=>	172,
		48084	=>	172,
		48085	=>	171,
		48086	=>	171,
		48087	=>	171,
		48088	=>	170,
		48089	=>	170,
		48090	=>	170,
		48091	=>	169,
		48092	=>	169,
		48093	=>	169,
		48094	=>	168,
		48095	=>	168,
		48096	=>	168,
		48097	=>	167,
		48098	=>	167,
		48099	=>	167,
		48100	=>	167,
		48101	=>	166,
		48102	=>	166,
		48103	=>	166,
		48104	=>	165,
		48105	=>	165,
		48106	=>	165,
		48107	=>	164,
		48108	=>	164,
		48109	=>	164,
		48110	=>	163,
		48111	=>	163,
		48112	=>	163,
		48113	=>	162,
		48114	=>	162,
		48115	=>	162,
		48116	=>	162,
		48117	=>	161,
		48118	=>	161,
		48119	=>	161,
		48120	=>	160,
		48121	=>	160,
		48122	=>	160,
		48123	=>	159,
		48124	=>	159,
		48125	=>	159,
		48126	=>	158,
		48127	=>	158,
		48128	=>	158,
		48129	=>	157,
		48130	=>	157,
		48131	=>	157,
		48132	=>	157,
		48133	=>	156,
		48134	=>	156,
		48135	=>	156,
		48136	=>	155,
		48137	=>	155,
		48138	=>	155,
		48139	=>	154,
		48140	=>	154,
		48141	=>	154,
		48142	=>	154,
		48143	=>	153,
		48144	=>	153,
		48145	=>	153,
		48146	=>	152,
		48147	=>	152,
		48148	=>	152,
		48149	=>	151,
		48150	=>	151,
		48151	=>	151,
		48152	=>	150,
		48153	=>	150,
		48154	=>	150,
		48155	=>	150,
		48156	=>	149,
		48157	=>	149,
		48158	=>	149,
		48159	=>	148,
		48160	=>	148,
		48161	=>	148,
		48162	=>	147,
		48163	=>	147,
		48164	=>	147,
		48165	=>	147,
		48166	=>	146,
		48167	=>	146,
		48168	=>	146,
		48169	=>	145,
		48170	=>	145,
		48171	=>	145,
		48172	=>	145,
		48173	=>	144,
		48174	=>	144,
		48175	=>	144,
		48176	=>	143,
		48177	=>	143,
		48178	=>	143,
		48179	=>	142,
		48180	=>	142,
		48181	=>	142,
		48182	=>	142,
		48183	=>	141,
		48184	=>	141,
		48185	=>	141,
		48186	=>	140,
		48187	=>	140,
		48188	=>	140,
		48189	=>	140,
		48190	=>	139,
		48191	=>	139,
		48192	=>	139,
		48193	=>	138,
		48194	=>	138,
		48195	=>	138,
		48196	=>	138,
		48197	=>	137,
		48198	=>	137,
		48199	=>	137,
		48200	=>	136,
		48201	=>	136,
		48202	=>	136,
		48203	=>	136,
		48204	=>	135,
		48205	=>	135,
		48206	=>	135,
		48207	=>	134,
		48208	=>	134,
		48209	=>	134,
		48210	=>	134,
		48211	=>	133,
		48212	=>	133,
		48213	=>	133,
		48214	=>	132,
		48215	=>	132,
		48216	=>	132,
		48217	=>	132,
		48218	=>	131,
		48219	=>	131,
		48220	=>	131,
		48221	=>	130,
		48222	=>	130,
		48223	=>	130,
		48224	=>	130,
		48225	=>	129,
		48226	=>	129,
		48227	=>	129,
		48228	=>	128,
		48229	=>	128,
		48230	=>	128,
		48231	=>	128,
		48232	=>	127,
		48233	=>	127,
		48234	=>	127,
		48235	=>	127,
		48236	=>	126,
		48237	=>	126,
		48238	=>	126,
		48239	=>	125,
		48240	=>	125,
		48241	=>	125,
		48242	=>	125,
		48243	=>	124,
		48244	=>	124,
		48245	=>	124,
		48246	=>	124,
		48247	=>	123,
		48248	=>	123,
		48249	=>	123,
		48250	=>	122,
		48251	=>	122,
		48252	=>	122,
		48253	=>	122,
		48254	=>	121,
		48255	=>	121,
		48256	=>	121,
		48257	=>	121,
		48258	=>	120,
		48259	=>	120,
		48260	=>	120,
		48261	=>	119,
		48262	=>	119,
		48263	=>	119,
		48264	=>	119,
		48265	=>	118,
		48266	=>	118,
		48267	=>	118,
		48268	=>	118,
		48269	=>	117,
		48270	=>	117,
		48271	=>	117,
		48272	=>	117,
		48273	=>	116,
		48274	=>	116,
		48275	=>	116,
		48276	=>	115,
		48277	=>	115,
		48278	=>	115,
		48279	=>	115,
		48280	=>	114,
		48281	=>	114,
		48282	=>	114,
		48283	=>	114,
		48284	=>	113,
		48285	=>	113,
		48286	=>	113,
		48287	=>	113,
		48288	=>	112,
		48289	=>	112,
		48290	=>	112,
		48291	=>	112,
		48292	=>	111,
		48293	=>	111,
		48294	=>	111,
		48295	=>	111,
		48296	=>	110,
		48297	=>	110,
		48298	=>	110,
		48299	=>	110,
		48300	=>	109,
		48301	=>	109,
		48302	=>	109,
		48303	=>	108,
		48304	=>	108,
		48305	=>	108,
		48306	=>	108,
		48307	=>	107,
		48308	=>	107,
		48309	=>	107,
		48310	=>	107,
		48311	=>	106,
		48312	=>	106,
		48313	=>	106,
		48314	=>	106,
		48315	=>	105,
		48316	=>	105,
		48317	=>	105,
		48318	=>	105,
		48319	=>	104,
		48320	=>	104,
		48321	=>	104,
		48322	=>	104,
		48323	=>	103,
		48324	=>	103,
		48325	=>	103,
		48326	=>	103,
		48327	=>	102,
		48328	=>	102,
		48329	=>	102,
		48330	=>	102,
		48331	=>	101,
		48332	=>	101,
		48333	=>	101,
		48334	=>	101,
		48335	=>	100,
		48336	=>	100,
		48337	=>	100,
		48338	=>	100,
		48339	=>	99,
		48340	=>	99,
		48341	=>	99,
		48342	=>	99,
		48343	=>	99,
		48344	=>	98,
		48345	=>	98,
		48346	=>	98,
		48347	=>	98,
		48348	=>	97,
		48349	=>	97,
		48350	=>	97,
		48351	=>	97,
		48352	=>	96,
		48353	=>	96,
		48354	=>	96,
		48355	=>	96,
		48356	=>	95,
		48357	=>	95,
		48358	=>	95,
		48359	=>	95,
		48360	=>	94,
		48361	=>	94,
		48362	=>	94,
		48363	=>	94,
		48364	=>	93,
		48365	=>	93,
		48366	=>	93,
		48367	=>	93,
		48368	=>	93,
		48369	=>	92,
		48370	=>	92,
		48371	=>	92,
		48372	=>	92,
		48373	=>	91,
		48374	=>	91,
		48375	=>	91,
		48376	=>	91,
		48377	=>	90,
		48378	=>	90,
		48379	=>	90,
		48380	=>	90,
		48381	=>	89,
		48382	=>	89,
		48383	=>	89,
		48384	=>	89,
		48385	=>	89,
		48386	=>	88,
		48387	=>	88,
		48388	=>	88,
		48389	=>	88,
		48390	=>	87,
		48391	=>	87,
		48392	=>	87,
		48393	=>	87,
		48394	=>	86,
		48395	=>	86,
		48396	=>	86,
		48397	=>	86,
		48398	=>	86,
		48399	=>	85,
		48400	=>	85,
		48401	=>	85,
		48402	=>	85,
		48403	=>	84,
		48404	=>	84,
		48405	=>	84,
		48406	=>	84,
		48407	=>	84,
		48408	=>	83,
		48409	=>	83,
		48410	=>	83,
		48411	=>	83,
		48412	=>	82,
		48413	=>	82,
		48414	=>	82,
		48415	=>	82,
		48416	=>	82,
		48417	=>	81,
		48418	=>	81,
		48419	=>	81,
		48420	=>	81,
		48421	=>	80,
		48422	=>	80,
		48423	=>	80,
		48424	=>	80,
		48425	=>	80,
		48426	=>	79,
		48427	=>	79,
		48428	=>	79,
		48429	=>	79,
		48430	=>	78,
		48431	=>	78,
		48432	=>	78,
		48433	=>	78,
		48434	=>	78,
		48435	=>	77,
		48436	=>	77,
		48437	=>	77,
		48438	=>	77,
		48439	=>	77,
		48440	=>	76,
		48441	=>	76,
		48442	=>	76,
		48443	=>	76,
		48444	=>	75,
		48445	=>	75,
		48446	=>	75,
		48447	=>	75,
		48448	=>	75,
		48449	=>	74,
		48450	=>	74,
		48451	=>	74,
		48452	=>	74,
		48453	=>	74,
		48454	=>	73,
		48455	=>	73,
		48456	=>	73,
		48457	=>	73,
		48458	=>	73,
		48459	=>	72,
		48460	=>	72,
		48461	=>	72,
		48462	=>	72,
		48463	=>	71,
		48464	=>	71,
		48465	=>	71,
		48466	=>	71,
		48467	=>	71,
		48468	=>	70,
		48469	=>	70,
		48470	=>	70,
		48471	=>	70,
		48472	=>	70,
		48473	=>	69,
		48474	=>	69,
		48475	=>	69,
		48476	=>	69,
		48477	=>	69,
		48478	=>	68,
		48479	=>	68,
		48480	=>	68,
		48481	=>	68,
		48482	=>	68,
		48483	=>	67,
		48484	=>	67,
		48485	=>	67,
		48486	=>	67,
		48487	=>	67,
		48488	=>	66,
		48489	=>	66,
		48490	=>	66,
		48491	=>	66,
		48492	=>	66,
		48493	=>	65,
		48494	=>	65,
		48495	=>	65,
		48496	=>	65,
		48497	=>	65,
		48498	=>	64,
		48499	=>	64,
		48500	=>	64,
		48501	=>	64,
		48502	=>	64,
		48503	=>	63,
		48504	=>	63,
		48505	=>	63,
		48506	=>	63,
		48507	=>	63,
		48508	=>	62,
		48509	=>	62,
		48510	=>	62,
		48511	=>	62,
		48512	=>	62,
		48513	=>	61,
		48514	=>	61,
		48515	=>	61,
		48516	=>	61,
		48517	=>	61,
		48518	=>	61,
		48519	=>	60,
		48520	=>	60,
		48521	=>	60,
		48522	=>	60,
		48523	=>	60,
		48524	=>	59,
		48525	=>	59,
		48526	=>	59,
		48527	=>	59,
		48528	=>	59,
		48529	=>	58,
		48530	=>	58,
		48531	=>	58,
		48532	=>	58,
		48533	=>	58,
		48534	=>	57,
		48535	=>	57,
		48536	=>	57,
		48537	=>	57,
		48538	=>	57,
		48539	=>	57,
		48540	=>	56,
		48541	=>	56,
		48542	=>	56,
		48543	=>	56,
		48544	=>	56,
		48545	=>	55,
		48546	=>	55,
		48547	=>	55,
		48548	=>	55,
		48549	=>	55,
		48550	=>	55,
		48551	=>	54,
		48552	=>	54,
		48553	=>	54,
		48554	=>	54,
		48555	=>	54,
		48556	=>	53,
		48557	=>	53,
		48558	=>	53,
		48559	=>	53,
		48560	=>	53,
		48561	=>	53,
		48562	=>	52,
		48563	=>	52,
		48564	=>	52,
		48565	=>	52,
		48566	=>	52,
		48567	=>	52,
		48568	=>	51,
		48569	=>	51,
		48570	=>	51,
		48571	=>	51,
		48572	=>	51,
		48573	=>	50,
		48574	=>	50,
		48575	=>	50,
		48576	=>	50,
		48577	=>	50,
		48578	=>	50,
		48579	=>	49,
		48580	=>	49,
		48581	=>	49,
		48582	=>	49,
		48583	=>	49,
		48584	=>	49,
		48585	=>	48,
		48586	=>	48,
		48587	=>	48,
		48588	=>	48,
		48589	=>	48,
		48590	=>	48,
		48591	=>	47,
		48592	=>	47,
		48593	=>	47,
		48594	=>	47,
		48595	=>	47,
		48596	=>	47,
		48597	=>	46,
		48598	=>	46,
		48599	=>	46,
		48600	=>	46,
		48601	=>	46,
		48602	=>	46,
		48603	=>	45,
		48604	=>	45,
		48605	=>	45,
		48606	=>	45,
		48607	=>	45,
		48608	=>	45,
		48609	=>	44,
		48610	=>	44,
		48611	=>	44,
		48612	=>	44,
		48613	=>	44,
		48614	=>	44,
		48615	=>	43,
		48616	=>	43,
		48617	=>	43,
		48618	=>	43,
		48619	=>	43,
		48620	=>	43,
		48621	=>	42,
		48622	=>	42,
		48623	=>	42,
		48624	=>	42,
		48625	=>	42,
		48626	=>	42,
		48627	=>	41,
		48628	=>	41,
		48629	=>	41,
		48630	=>	41,
		48631	=>	41,
		48632	=>	41,
		48633	=>	41,
		48634	=>	40,
		48635	=>	40,
		48636	=>	40,
		48637	=>	40,
		48638	=>	40,
		48639	=>	40,
		48640	=>	39,
		48641	=>	39,
		48642	=>	39,
		48643	=>	39,
		48644	=>	39,
		48645	=>	39,
		48646	=>	39,
		48647	=>	38,
		48648	=>	38,
		48649	=>	38,
		48650	=>	38,
		48651	=>	38,
		48652	=>	38,
		48653	=>	37,
		48654	=>	37,
		48655	=>	37,
		48656	=>	37,
		48657	=>	37,
		48658	=>	37,
		48659	=>	37,
		48660	=>	36,
		48661	=>	36,
		48662	=>	36,
		48663	=>	36,
		48664	=>	36,
		48665	=>	36,
		48666	=>	36,
		48667	=>	35,
		48668	=>	35,
		48669	=>	35,
		48670	=>	35,
		48671	=>	35,
		48672	=>	35,
		48673	=>	35,
		48674	=>	34,
		48675	=>	34,
		48676	=>	34,
		48677	=>	34,
		48678	=>	34,
		48679	=>	34,
		48680	=>	34,
		48681	=>	33,
		48682	=>	33,
		48683	=>	33,
		48684	=>	33,
		48685	=>	33,
		48686	=>	33,
		48687	=>	33,
		48688	=>	32,
		48689	=>	32,
		48690	=>	32,
		48691	=>	32,
		48692	=>	32,
		48693	=>	32,
		48694	=>	32,
		48695	=>	31,
		48696	=>	31,
		48697	=>	31,
		48698	=>	31,
		48699	=>	31,
		48700	=>	31,
		48701	=>	31,
		48702	=>	30,
		48703	=>	30,
		48704	=>	30,
		48705	=>	30,
		48706	=>	30,
		48707	=>	30,
		48708	=>	30,
		48709	=>	30,
		48710	=>	29,
		48711	=>	29,
		48712	=>	29,
		48713	=>	29,
		48714	=>	29,
		48715	=>	29,
		48716	=>	29,
		48717	=>	28,
		48718	=>	28,
		48719	=>	28,
		48720	=>	28,
		48721	=>	28,
		48722	=>	28,
		48723	=>	28,
		48724	=>	28,
		48725	=>	27,
		48726	=>	27,
		48727	=>	27,
		48728	=>	27,
		48729	=>	27,
		48730	=>	27,
		48731	=>	27,
		48732	=>	27,
		48733	=>	26,
		48734	=>	26,
		48735	=>	26,
		48736	=>	26,
		48737	=>	26,
		48738	=>	26,
		48739	=>	26,
		48740	=>	26,
		48741	=>	25,
		48742	=>	25,
		48743	=>	25,
		48744	=>	25,
		48745	=>	25,
		48746	=>	25,
		48747	=>	25,
		48748	=>	25,
		48749	=>	24,
		48750	=>	24,
		48751	=>	24,
		48752	=>	24,
		48753	=>	24,
		48754	=>	24,
		48755	=>	24,
		48756	=>	24,
		48757	=>	23,
		48758	=>	23,
		48759	=>	23,
		48760	=>	23,
		48761	=>	23,
		48762	=>	23,
		48763	=>	23,
		48764	=>	23,
		48765	=>	23,
		48766	=>	22,
		48767	=>	22,
		48768	=>	22,
		48769	=>	22,
		48770	=>	22,
		48771	=>	22,
		48772	=>	22,
		48773	=>	22,
		48774	=>	22,
		48775	=>	21,
		48776	=>	21,
		48777	=>	21,
		48778	=>	21,
		48779	=>	21,
		48780	=>	21,
		48781	=>	21,
		48782	=>	21,
		48783	=>	21,
		48784	=>	20,
		48785	=>	20,
		48786	=>	20,
		48787	=>	20,
		48788	=>	20,
		48789	=>	20,
		48790	=>	20,
		48791	=>	20,
		48792	=>	20,
		48793	=>	19,
		48794	=>	19,
		48795	=>	19,
		48796	=>	19,
		48797	=>	19,
		48798	=>	19,
		48799	=>	19,
		48800	=>	19,
		48801	=>	19,
		48802	=>	18,
		48803	=>	18,
		48804	=>	18,
		48805	=>	18,
		48806	=>	18,
		48807	=>	18,
		48808	=>	18,
		48809	=>	18,
		48810	=>	18,
		48811	=>	18,
		48812	=>	17,
		48813	=>	17,
		48814	=>	17,
		48815	=>	17,
		48816	=>	17,
		48817	=>	17,
		48818	=>	17,
		48819	=>	17,
		48820	=>	17,
		48821	=>	16,
		48822	=>	16,
		48823	=>	16,
		48824	=>	16,
		48825	=>	16,
		48826	=>	16,
		48827	=>	16,
		48828	=>	16,
		48829	=>	16,
		48830	=>	16,
		48831	=>	16,
		48832	=>	15,
		48833	=>	15,
		48834	=>	15,
		48835	=>	15,
		48836	=>	15,
		48837	=>	15,
		48838	=>	15,
		48839	=>	15,
		48840	=>	15,
		48841	=>	15,
		48842	=>	14,
		48843	=>	14,
		48844	=>	14,
		48845	=>	14,
		48846	=>	14,
		48847	=>	14,
		48848	=>	14,
		48849	=>	14,
		48850	=>	14,
		48851	=>	14,
		48852	=>	14,
		48853	=>	13,
		48854	=>	13,
		48855	=>	13,
		48856	=>	13,
		48857	=>	13,
		48858	=>	13,
		48859	=>	13,
		48860	=>	13,
		48861	=>	13,
		48862	=>	13,
		48863	=>	13,
		48864	=>	12,
		48865	=>	12,
		48866	=>	12,
		48867	=>	12,
		48868	=>	12,
		48869	=>	12,
		48870	=>	12,
		48871	=>	12,
		48872	=>	12,
		48873	=>	12,
		48874	=>	12,
		48875	=>	12,
		48876	=>	11,
		48877	=>	11,
		48878	=>	11,
		48879	=>	11,
		48880	=>	11,
		48881	=>	11,
		48882	=>	11,
		48883	=>	11,
		48884	=>	11,
		48885	=>	11,
		48886	=>	11,
		48887	=>	11,
		48888	=>	10,
		48889	=>	10,
		48890	=>	10,
		48891	=>	10,
		48892	=>	10,
		48893	=>	10,
		48894	=>	10,
		48895	=>	10,
		48896	=>	10,
		48897	=>	10,
		48898	=>	10,
		48899	=>	10,
		48900	=>	10,
		48901	=>	9,
		48902	=>	9,
		48903	=>	9,
		48904	=>	9,
		48905	=>	9,
		48906	=>	9,
		48907	=>	9,
		48908	=>	9,
		48909	=>	9,
		48910	=>	9,
		48911	=>	9,
		48912	=>	9,
		48913	=>	9,
		48914	=>	9,
		48915	=>	8,
		48916	=>	8,
		48917	=>	8,
		48918	=>	8,
		48919	=>	8,
		48920	=>	8,
		48921	=>	8,
		48922	=>	8,
		48923	=>	8,
		48924	=>	8,
		48925	=>	8,
		48926	=>	8,
		48927	=>	8,
		48928	=>	8,
		48929	=>	7,
		48930	=>	7,
		48931	=>	7,
		48932	=>	7,
		48933	=>	7,
		48934	=>	7,
		48935	=>	7,
		48936	=>	7,
		48937	=>	7,
		48938	=>	7,
		48939	=>	7,
		48940	=>	7,
		48941	=>	7,
		48942	=>	7,
		48943	=>	7,
		48944	=>	7,
		48945	=>	6,
		48946	=>	6,
		48947	=>	6,
		48948	=>	6,
		48949	=>	6,
		48950	=>	6,
		48951	=>	6,
		48952	=>	6,
		48953	=>	6,
		48954	=>	6,
		48955	=>	6,
		48956	=>	6,
		48957	=>	6,
		48958	=>	6,
		48959	=>	6,
		48960	=>	6,
		48961	=>	5,
		48962	=>	5,
		48963	=>	5,
		48964	=>	5,
		48965	=>	5,
		48966	=>	5,
		48967	=>	5,
		48968	=>	5,
		48969	=>	5,
		48970	=>	5,
		48971	=>	5,
		48972	=>	5,
		48973	=>	5,
		48974	=>	5,
		48975	=>	5,
		48976	=>	5,
		48977	=>	5,
		48978	=>	5,
		48979	=>	5,
		48980	=>	4,
		48981	=>	4,
		48982	=>	4,
		48983	=>	4,
		48984	=>	4,
		48985	=>	4,
		48986	=>	4,
		48987	=>	4,
		48988	=>	4,
		48989	=>	4,
		48990	=>	4,
		48991	=>	4,
		48992	=>	4,
		48993	=>	4,
		48994	=>	4,
		48995	=>	4,
		48996	=>	4,
		48997	=>	4,
		48998	=>	4,
		48999	=>	4,
		49000	=>	3,
		49001	=>	3,
		49002	=>	3,
		49003	=>	3,
		49004	=>	3,
		49005	=>	3,
		49006	=>	3,
		49007	=>	3,
		49008	=>	3,
		49009	=>	3,
		49010	=>	3,
		49011	=>	3,
		49012	=>	3,
		49013	=>	3,
		49014	=>	3,
		49015	=>	3,
		49016	=>	3,
		49017	=>	3,
		49018	=>	3,
		49019	=>	3,
		49020	=>	3,
		49021	=>	3,
		49022	=>	3,
		49023	=>	3,
		49024	=>	2,
		49025	=>	2,
		49026	=>	2,
		49027	=>	2,
		49028	=>	2,
		49029	=>	2,
		49030	=>	2,
		49031	=>	2,
		49032	=>	2,
		49033	=>	2,
		49034	=>	2,
		49035	=>	2,
		49036	=>	2,
		49037	=>	2,
		49038	=>	2,
		49039	=>	2,
		49040	=>	2,
		49041	=>	2,
		49042	=>	2,
		49043	=>	2,
		49044	=>	2,
		49045	=>	2,
		49046	=>	2,
		49047	=>	2,
		49048	=>	2,
		49049	=>	2,
		49050	=>	2,
		49051	=>	2,
		49052	=>	2,
		49053	=>	1,
		49054	=>	1,
		49055	=>	1,
		49056	=>	1,
		49057	=>	1,
		49058	=>	1,
		49059	=>	1,
		49060	=>	1,
		49061	=>	1,
		49062	=>	1,
		49063	=>	1,
		49064	=>	1,
		49065	=>	1,
		49066	=>	1,
		49067	=>	1,
		49068	=>	1,
		49069	=>	1,
		49070	=>	1,
		49071	=>	1,
		49072	=>	1,
		49073	=>	1,
		49074	=>	1,
		49075	=>	1,
		49076	=>	1,
		49077	=>	1,
		49078	=>	1,
		49079	=>	1,
		49080	=>	1,
		49081	=>	1,
		49082	=>	1,
		49083	=>	1,
		49084	=>	1,
		49085	=>	1,
		49086	=>	1,
		49087	=>	1,
		49088	=>	1,
		49089	=>	1,
		49090	=>	1,
		49091	=>	1,
		49092	=>	1,
		49093	=>	1,
		49094	=>	1,
		49095	=>	0,
		49096	=>	0,
		49097	=>	0,
		49098	=>	0,
		49099	=>	0,
		49100	=>	0,
		49101	=>	0,
		49102	=>	0,
		49103	=>	0,
		49104	=>	0,
		49105	=>	0,
		49106	=>	0,
		49107	=>	0,
		49108	=>	0,
		49109	=>	0,
		49110	=>	0,
		49111	=>	0,
		49112	=>	0,
		49113	=>	0,
		49114	=>	0,
		49115	=>	0,
		49116	=>	0,
		49117	=>	0,
		49118	=>	0,
		49119	=>	0,
		49120	=>	0,
		49121	=>	0,
		49122	=>	0,
		49123	=>	0,
		49124	=>	0,
		49125	=>	0,
		49126	=>	0,
		49127	=>	0,
		49128	=>	0,
		49129	=>	0,
		49130	=>	0,
		49131	=>	0,
		49132	=>	0,
		49133	=>	0,
		49134	=>	0,
		49135	=>	0,
		49136	=>	0,
		49137	=>	0,
		49138	=>	0,
		49139	=>	0,
		49140	=>	0,
		49141	=>	0,
		49142	=>	0,
		49143	=>	0,
		49144	=>	0,
		49145	=>	0,
		49146	=>	0,
		49147	=>	0,
		49148	=>	0,
		49149	=>	0,
		49150	=>	0,
		49151	=>	0,
		49152	=>	0,
		49153	=>	0,
		49154	=>	0,
		49155	=>	0,
		49156	=>	0,
		49157	=>	0,
		49158	=>	0,
		49159	=>	0,
		49160	=>	0,
		49161	=>	0,
		49162	=>	0,
		49163	=>	0,
		49164	=>	0,
		49165	=>	0,
		49166	=>	0,
		49167	=>	0,
		49168	=>	0,
		49169	=>	0,
		49170	=>	0,
		49171	=>	0,
		49172	=>	0,
		49173	=>	0,
		49174	=>	0,
		49175	=>	0,
		49176	=>	0,
		49177	=>	0,
		49178	=>	0,
		49179	=>	0,
		49180	=>	0,
		49181	=>	0,
		49182	=>	0,
		49183	=>	0,
		49184	=>	0,
		49185	=>	0,
		49186	=>	0,
		49187	=>	0,
		49188	=>	0,
		49189	=>	0,
		49190	=>	0,
		49191	=>	0,
		49192	=>	0,
		49193	=>	0,
		49194	=>	0,
		49195	=>	0,
		49196	=>	0,
		49197	=>	0,
		49198	=>	0,
		49199	=>	0,
		49200	=>	0,
		49201	=>	0,
		49202	=>	0,
		49203	=>	0,
		49204	=>	0,
		49205	=>	0,
		49206	=>	0,
		49207	=>	0,
		49208	=>	0,
		49209	=>	0,
		49210	=>	1,
		49211	=>	1,
		49212	=>	1,
		49213	=>	1,
		49214	=>	1,
		49215	=>	1,
		49216	=>	1,
		49217	=>	1,
		49218	=>	1,
		49219	=>	1,
		49220	=>	1,
		49221	=>	1,
		49222	=>	1,
		49223	=>	1,
		49224	=>	1,
		49225	=>	1,
		49226	=>	1,
		49227	=>	1,
		49228	=>	1,
		49229	=>	1,
		49230	=>	1,
		49231	=>	1,
		49232	=>	1,
		49233	=>	1,
		49234	=>	1,
		49235	=>	1,
		49236	=>	1,
		49237	=>	1,
		49238	=>	1,
		49239	=>	1,
		49240	=>	1,
		49241	=>	1,
		49242	=>	1,
		49243	=>	1,
		49244	=>	1,
		49245	=>	1,
		49246	=>	1,
		49247	=>	1,
		49248	=>	1,
		49249	=>	1,
		49250	=>	1,
		49251	=>	1,
		49252	=>	2,
		49253	=>	2,
		49254	=>	2,
		49255	=>	2,
		49256	=>	2,
		49257	=>	2,
		49258	=>	2,
		49259	=>	2,
		49260	=>	2,
		49261	=>	2,
		49262	=>	2,
		49263	=>	2,
		49264	=>	2,
		49265	=>	2,
		49266	=>	2,
		49267	=>	2,
		49268	=>	2,
		49269	=>	2,
		49270	=>	2,
		49271	=>	2,
		49272	=>	2,
		49273	=>	2,
		49274	=>	2,
		49275	=>	2,
		49276	=>	2,
		49277	=>	2,
		49278	=>	2,
		49279	=>	2,
		49280	=>	2,
		49281	=>	3,
		49282	=>	3,
		49283	=>	3,
		49284	=>	3,
		49285	=>	3,
		49286	=>	3,
		49287	=>	3,
		49288	=>	3,
		49289	=>	3,
		49290	=>	3,
		49291	=>	3,
		49292	=>	3,
		49293	=>	3,
		49294	=>	3,
		49295	=>	3,
		49296	=>	3,
		49297	=>	3,
		49298	=>	3,
		49299	=>	3,
		49300	=>	3,
		49301	=>	3,
		49302	=>	3,
		49303	=>	3,
		49304	=>	3,
		49305	=>	4,
		49306	=>	4,
		49307	=>	4,
		49308	=>	4,
		49309	=>	4,
		49310	=>	4,
		49311	=>	4,
		49312	=>	4,
		49313	=>	4,
		49314	=>	4,
		49315	=>	4,
		49316	=>	4,
		49317	=>	4,
		49318	=>	4,
		49319	=>	4,
		49320	=>	4,
		49321	=>	4,
		49322	=>	4,
		49323	=>	4,
		49324	=>	4,
		49325	=>	5,
		49326	=>	5,
		49327	=>	5,
		49328	=>	5,
		49329	=>	5,
		49330	=>	5,
		49331	=>	5,
		49332	=>	5,
		49333	=>	5,
		49334	=>	5,
		49335	=>	5,
		49336	=>	5,
		49337	=>	5,
		49338	=>	5,
		49339	=>	5,
		49340	=>	5,
		49341	=>	5,
		49342	=>	5,
		49343	=>	5,
		49344	=>	6,
		49345	=>	6,
		49346	=>	6,
		49347	=>	6,
		49348	=>	6,
		49349	=>	6,
		49350	=>	6,
		49351	=>	6,
		49352	=>	6,
		49353	=>	6,
		49354	=>	6,
		49355	=>	6,
		49356	=>	6,
		49357	=>	6,
		49358	=>	6,
		49359	=>	6,
		49360	=>	7,
		49361	=>	7,
		49362	=>	7,
		49363	=>	7,
		49364	=>	7,
		49365	=>	7,
		49366	=>	7,
		49367	=>	7,
		49368	=>	7,
		49369	=>	7,
		49370	=>	7,
		49371	=>	7,
		49372	=>	7,
		49373	=>	7,
		49374	=>	7,
		49375	=>	7,
		49376	=>	8,
		49377	=>	8,
		49378	=>	8,
		49379	=>	8,
		49380	=>	8,
		49381	=>	8,
		49382	=>	8,
		49383	=>	8,
		49384	=>	8,
		49385	=>	8,
		49386	=>	8,
		49387	=>	8,
		49388	=>	8,
		49389	=>	8,
		49390	=>	9,
		49391	=>	9,
		49392	=>	9,
		49393	=>	9,
		49394	=>	9,
		49395	=>	9,
		49396	=>	9,
		49397	=>	9,
		49398	=>	9,
		49399	=>	9,
		49400	=>	9,
		49401	=>	9,
		49402	=>	9,
		49403	=>	9,
		49404	=>	10,
		49405	=>	10,
		49406	=>	10,
		49407	=>	10,
		49408	=>	10,
		49409	=>	10,
		49410	=>	10,
		49411	=>	10,
		49412	=>	10,
		49413	=>	10,
		49414	=>	10,
		49415	=>	10,
		49416	=>	10,
		49417	=>	11,
		49418	=>	11,
		49419	=>	11,
		49420	=>	11,
		49421	=>	11,
		49422	=>	11,
		49423	=>	11,
		49424	=>	11,
		49425	=>	11,
		49426	=>	11,
		49427	=>	11,
		49428	=>	11,
		49429	=>	12,
		49430	=>	12,
		49431	=>	12,
		49432	=>	12,
		49433	=>	12,
		49434	=>	12,
		49435	=>	12,
		49436	=>	12,
		49437	=>	12,
		49438	=>	12,
		49439	=>	12,
		49440	=>	12,
		49441	=>	13,
		49442	=>	13,
		49443	=>	13,
		49444	=>	13,
		49445	=>	13,
		49446	=>	13,
		49447	=>	13,
		49448	=>	13,
		49449	=>	13,
		49450	=>	13,
		49451	=>	13,
		49452	=>	14,
		49453	=>	14,
		49454	=>	14,
		49455	=>	14,
		49456	=>	14,
		49457	=>	14,
		49458	=>	14,
		49459	=>	14,
		49460	=>	14,
		49461	=>	14,
		49462	=>	14,
		49463	=>	15,
		49464	=>	15,
		49465	=>	15,
		49466	=>	15,
		49467	=>	15,
		49468	=>	15,
		49469	=>	15,
		49470	=>	15,
		49471	=>	15,
		49472	=>	15,
		49473	=>	16,
		49474	=>	16,
		49475	=>	16,
		49476	=>	16,
		49477	=>	16,
		49478	=>	16,
		49479	=>	16,
		49480	=>	16,
		49481	=>	16,
		49482	=>	16,
		49483	=>	16,
		49484	=>	17,
		49485	=>	17,
		49486	=>	17,
		49487	=>	17,
		49488	=>	17,
		49489	=>	17,
		49490	=>	17,
		49491	=>	17,
		49492	=>	17,
		49493	=>	18,
		49494	=>	18,
		49495	=>	18,
		49496	=>	18,
		49497	=>	18,
		49498	=>	18,
		49499	=>	18,
		49500	=>	18,
		49501	=>	18,
		49502	=>	18,
		49503	=>	19,
		49504	=>	19,
		49505	=>	19,
		49506	=>	19,
		49507	=>	19,
		49508	=>	19,
		49509	=>	19,
		49510	=>	19,
		49511	=>	19,
		49512	=>	20,
		49513	=>	20,
		49514	=>	20,
		49515	=>	20,
		49516	=>	20,
		49517	=>	20,
		49518	=>	20,
		49519	=>	20,
		49520	=>	20,
		49521	=>	21,
		49522	=>	21,
		49523	=>	21,
		49524	=>	21,
		49525	=>	21,
		49526	=>	21,
		49527	=>	21,
		49528	=>	21,
		49529	=>	21,
		49530	=>	22,
		49531	=>	22,
		49532	=>	22,
		49533	=>	22,
		49534	=>	22,
		49535	=>	22,
		49536	=>	22,
		49537	=>	22,
		49538	=>	22,
		49539	=>	23,
		49540	=>	23,
		49541	=>	23,
		49542	=>	23,
		49543	=>	23,
		49544	=>	23,
		49545	=>	23,
		49546	=>	23,
		49547	=>	23,
		49548	=>	24,
		49549	=>	24,
		49550	=>	24,
		49551	=>	24,
		49552	=>	24,
		49553	=>	24,
		49554	=>	24,
		49555	=>	24,
		49556	=>	25,
		49557	=>	25,
		49558	=>	25,
		49559	=>	25,
		49560	=>	25,
		49561	=>	25,
		49562	=>	25,
		49563	=>	25,
		49564	=>	26,
		49565	=>	26,
		49566	=>	26,
		49567	=>	26,
		49568	=>	26,
		49569	=>	26,
		49570	=>	26,
		49571	=>	26,
		49572	=>	27,
		49573	=>	27,
		49574	=>	27,
		49575	=>	27,
		49576	=>	27,
		49577	=>	27,
		49578	=>	27,
		49579	=>	27,
		49580	=>	28,
		49581	=>	28,
		49582	=>	28,
		49583	=>	28,
		49584	=>	28,
		49585	=>	28,
		49586	=>	28,
		49587	=>	28,
		49588	=>	29,
		49589	=>	29,
		49590	=>	29,
		49591	=>	29,
		49592	=>	29,
		49593	=>	29,
		49594	=>	29,
		49595	=>	30,
		49596	=>	30,
		49597	=>	30,
		49598	=>	30,
		49599	=>	30,
		49600	=>	30,
		49601	=>	30,
		49602	=>	30,
		49603	=>	31,
		49604	=>	31,
		49605	=>	31,
		49606	=>	31,
		49607	=>	31,
		49608	=>	31,
		49609	=>	31,
		49610	=>	32,
		49611	=>	32,
		49612	=>	32,
		49613	=>	32,
		49614	=>	32,
		49615	=>	32,
		49616	=>	32,
		49617	=>	33,
		49618	=>	33,
		49619	=>	33,
		49620	=>	33,
		49621	=>	33,
		49622	=>	33,
		49623	=>	33,
		49624	=>	34,
		49625	=>	34,
		49626	=>	34,
		49627	=>	34,
		49628	=>	34,
		49629	=>	34,
		49630	=>	34,
		49631	=>	35,
		49632	=>	35,
		49633	=>	35,
		49634	=>	35,
		49635	=>	35,
		49636	=>	35,
		49637	=>	35,
		49638	=>	36,
		49639	=>	36,
		49640	=>	36,
		49641	=>	36,
		49642	=>	36,
		49643	=>	36,
		49644	=>	36,
		49645	=>	37,
		49646	=>	37,
		49647	=>	37,
		49648	=>	37,
		49649	=>	37,
		49650	=>	37,
		49651	=>	37,
		49652	=>	38,
		49653	=>	38,
		49654	=>	38,
		49655	=>	38,
		49656	=>	38,
		49657	=>	38,
		49658	=>	39,
		49659	=>	39,
		49660	=>	39,
		49661	=>	39,
		49662	=>	39,
		49663	=>	39,
		49664	=>	39,
		49665	=>	40,
		49666	=>	40,
		49667	=>	40,
		49668	=>	40,
		49669	=>	40,
		49670	=>	40,
		49671	=>	41,
		49672	=>	41,
		49673	=>	41,
		49674	=>	41,
		49675	=>	41,
		49676	=>	41,
		49677	=>	41,
		49678	=>	42,
		49679	=>	42,
		49680	=>	42,
		49681	=>	42,
		49682	=>	42,
		49683	=>	42,
		49684	=>	43,
		49685	=>	43,
		49686	=>	43,
		49687	=>	43,
		49688	=>	43,
		49689	=>	43,
		49690	=>	44,
		49691	=>	44,
		49692	=>	44,
		49693	=>	44,
		49694	=>	44,
		49695	=>	44,
		49696	=>	45,
		49697	=>	45,
		49698	=>	45,
		49699	=>	45,
		49700	=>	45,
		49701	=>	45,
		49702	=>	46,
		49703	=>	46,
		49704	=>	46,
		49705	=>	46,
		49706	=>	46,
		49707	=>	46,
		49708	=>	47,
		49709	=>	47,
		49710	=>	47,
		49711	=>	47,
		49712	=>	47,
		49713	=>	47,
		49714	=>	48,
		49715	=>	48,
		49716	=>	48,
		49717	=>	48,
		49718	=>	48,
		49719	=>	48,
		49720	=>	49,
		49721	=>	49,
		49722	=>	49,
		49723	=>	49,
		49724	=>	49,
		49725	=>	49,
		49726	=>	50,
		49727	=>	50,
		49728	=>	50,
		49729	=>	50,
		49730	=>	50,
		49731	=>	50,
		49732	=>	51,
		49733	=>	51,
		49734	=>	51,
		49735	=>	51,
		49736	=>	51,
		49737	=>	52,
		49738	=>	52,
		49739	=>	52,
		49740	=>	52,
		49741	=>	52,
		49742	=>	52,
		49743	=>	53,
		49744	=>	53,
		49745	=>	53,
		49746	=>	53,
		49747	=>	53,
		49748	=>	53,
		49749	=>	54,
		49750	=>	54,
		49751	=>	54,
		49752	=>	54,
		49753	=>	54,
		49754	=>	55,
		49755	=>	55,
		49756	=>	55,
		49757	=>	55,
		49758	=>	55,
		49759	=>	55,
		49760	=>	56,
		49761	=>	56,
		49762	=>	56,
		49763	=>	56,
		49764	=>	56,
		49765	=>	57,
		49766	=>	57,
		49767	=>	57,
		49768	=>	57,
		49769	=>	57,
		49770	=>	57,
		49771	=>	58,
		49772	=>	58,
		49773	=>	58,
		49774	=>	58,
		49775	=>	58,
		49776	=>	59,
		49777	=>	59,
		49778	=>	59,
		49779	=>	59,
		49780	=>	59,
		49781	=>	60,
		49782	=>	60,
		49783	=>	60,
		49784	=>	60,
		49785	=>	60,
		49786	=>	61,
		49787	=>	61,
		49788	=>	61,
		49789	=>	61,
		49790	=>	61,
		49791	=>	61,
		49792	=>	62,
		49793	=>	62,
		49794	=>	62,
		49795	=>	62,
		49796	=>	62,
		49797	=>	63,
		49798	=>	63,
		49799	=>	63,
		49800	=>	63,
		49801	=>	63,
		49802	=>	64,
		49803	=>	64,
		49804	=>	64,
		49805	=>	64,
		49806	=>	64,
		49807	=>	65,
		49808	=>	65,
		49809	=>	65,
		49810	=>	65,
		49811	=>	65,
		49812	=>	66,
		49813	=>	66,
		49814	=>	66,
		49815	=>	66,
		49816	=>	66,
		49817	=>	67,
		49818	=>	67,
		49819	=>	67,
		49820	=>	67,
		49821	=>	67,
		49822	=>	68,
		49823	=>	68,
		49824	=>	68,
		49825	=>	68,
		49826	=>	68,
		49827	=>	69,
		49828	=>	69,
		49829	=>	69,
		49830	=>	69,
		49831	=>	69,
		49832	=>	70,
		49833	=>	70,
		49834	=>	70,
		49835	=>	70,
		49836	=>	70,
		49837	=>	71,
		49838	=>	71,
		49839	=>	71,
		49840	=>	71,
		49841	=>	71,
		49842	=>	72,
		49843	=>	72,
		49844	=>	72,
		49845	=>	72,
		49846	=>	73,
		49847	=>	73,
		49848	=>	73,
		49849	=>	73,
		49850	=>	73,
		49851	=>	74,
		49852	=>	74,
		49853	=>	74,
		49854	=>	74,
		49855	=>	74,
		49856	=>	75,
		49857	=>	75,
		49858	=>	75,
		49859	=>	75,
		49860	=>	75,
		49861	=>	76,
		49862	=>	76,
		49863	=>	76,
		49864	=>	76,
		49865	=>	77,
		49866	=>	77,
		49867	=>	77,
		49868	=>	77,
		49869	=>	77,
		49870	=>	78,
		49871	=>	78,
		49872	=>	78,
		49873	=>	78,
		49874	=>	78,
		49875	=>	79,
		49876	=>	79,
		49877	=>	79,
		49878	=>	79,
		49879	=>	80,
		49880	=>	80,
		49881	=>	80,
		49882	=>	80,
		49883	=>	80,
		49884	=>	81,
		49885	=>	81,
		49886	=>	81,
		49887	=>	81,
		49888	=>	82,
		49889	=>	82,
		49890	=>	82,
		49891	=>	82,
		49892	=>	82,
		49893	=>	83,
		49894	=>	83,
		49895	=>	83,
		49896	=>	83,
		49897	=>	84,
		49898	=>	84,
		49899	=>	84,
		49900	=>	84,
		49901	=>	84,
		49902	=>	85,
		49903	=>	85,
		49904	=>	85,
		49905	=>	85,
		49906	=>	86,
		49907	=>	86,
		49908	=>	86,
		49909	=>	86,
		49910	=>	86,
		49911	=>	87,
		49912	=>	87,
		49913	=>	87,
		49914	=>	87,
		49915	=>	88,
		49916	=>	88,
		49917	=>	88,
		49918	=>	88,
		49919	=>	89,
		49920	=>	89,
		49921	=>	89,
		49922	=>	89,
		49923	=>	89,
		49924	=>	90,
		49925	=>	90,
		49926	=>	90,
		49927	=>	90,
		49928	=>	91,
		49929	=>	91,
		49930	=>	91,
		49931	=>	91,
		49932	=>	92,
		49933	=>	92,
		49934	=>	92,
		49935	=>	92,
		49936	=>	93,
		49937	=>	93,
		49938	=>	93,
		49939	=>	93,
		49940	=>	93,
		49941	=>	94,
		49942	=>	94,
		49943	=>	94,
		49944	=>	94,
		49945	=>	95,
		49946	=>	95,
		49947	=>	95,
		49948	=>	95,
		49949	=>	96,
		49950	=>	96,
		49951	=>	96,
		49952	=>	96,
		49953	=>	97,
		49954	=>	97,
		49955	=>	97,
		49956	=>	97,
		49957	=>	98,
		49958	=>	98,
		49959	=>	98,
		49960	=>	98,
		49961	=>	99,
		49962	=>	99,
		49963	=>	99,
		49964	=>	99,
		49965	=>	99,
		49966	=>	100,
		49967	=>	100,
		49968	=>	100,
		49969	=>	100,
		49970	=>	101,
		49971	=>	101,
		49972	=>	101,
		49973	=>	101,
		49974	=>	102,
		49975	=>	102,
		49976	=>	102,
		49977	=>	102,
		49978	=>	103,
		49979	=>	103,
		49980	=>	103,
		49981	=>	103,
		49982	=>	104,
		49983	=>	104,
		49984	=>	104,
		49985	=>	104,
		49986	=>	105,
		49987	=>	105,
		49988	=>	105,
		49989	=>	105,
		49990	=>	106,
		49991	=>	106,
		49992	=>	106,
		49993	=>	106,
		49994	=>	107,
		49995	=>	107,
		49996	=>	107,
		49997	=>	107,
		49998	=>	108,
		49999	=>	108,
		50000	=>	108,
		50001	=>	108,
		50002	=>	109,
		50003	=>	109,
		50004	=>	109,
		50005	=>	110,
		50006	=>	110,
		50007	=>	110,
		50008	=>	110,
		50009	=>	111,
		50010	=>	111,
		50011	=>	111,
		50012	=>	111,
		50013	=>	112,
		50014	=>	112,
		50015	=>	112,
		50016	=>	112,
		50017	=>	113,
		50018	=>	113,
		50019	=>	113,
		50020	=>	113,
		50021	=>	114,
		50022	=>	114,
		50023	=>	114,
		50024	=>	114,
		50025	=>	115,
		50026	=>	115,
		50027	=>	115,
		50028	=>	115,
		50029	=>	116,
		50030	=>	116,
		50031	=>	116,
		50032	=>	117,
		50033	=>	117,
		50034	=>	117,
		50035	=>	117,
		50036	=>	118,
		50037	=>	118,
		50038	=>	118,
		50039	=>	118,
		50040	=>	119,
		50041	=>	119,
		50042	=>	119,
		50043	=>	119,
		50044	=>	120,
		50045	=>	120,
		50046	=>	120,
		50047	=>	121,
		50048	=>	121,
		50049	=>	121,
		50050	=>	121,
		50051	=>	122,
		50052	=>	122,
		50053	=>	122,
		50054	=>	122,
		50055	=>	123,
		50056	=>	123,
		50057	=>	123,
		50058	=>	124,
		50059	=>	124,
		50060	=>	124,
		50061	=>	124,
		50062	=>	125,
		50063	=>	125,
		50064	=>	125,
		50065	=>	125,
		50066	=>	126,
		50067	=>	126,
		50068	=>	126,
		50069	=>	127,
		50070	=>	127,
		50071	=>	127,
		50072	=>	127,
		50073	=>	128,
		50074	=>	128,
		50075	=>	128,
		50076	=>	128,
		50077	=>	129,
		50078	=>	129,
		50079	=>	129,
		50080	=>	130,
		50081	=>	130,
		50082	=>	130,
		50083	=>	130,
		50084	=>	131,
		50085	=>	131,
		50086	=>	131,
		50087	=>	132,
		50088	=>	132,
		50089	=>	132,
		50090	=>	132,
		50091	=>	133,
		50092	=>	133,
		50093	=>	133,
		50094	=>	134,
		50095	=>	134,
		50096	=>	134,
		50097	=>	134,
		50098	=>	135,
		50099	=>	135,
		50100	=>	135,
		50101	=>	136,
		50102	=>	136,
		50103	=>	136,
		50104	=>	136,
		50105	=>	137,
		50106	=>	137,
		50107	=>	137,
		50108	=>	138,
		50109	=>	138,
		50110	=>	138,
		50111	=>	138,
		50112	=>	139,
		50113	=>	139,
		50114	=>	139,
		50115	=>	140,
		50116	=>	140,
		50117	=>	140,
		50118	=>	140,
		50119	=>	141,
		50120	=>	141,
		50121	=>	141,
		50122	=>	142,
		50123	=>	142,
		50124	=>	142,
		50125	=>	142,
		50126	=>	143,
		50127	=>	143,
		50128	=>	143,
		50129	=>	144,
		50130	=>	144,
		50131	=>	144,
		50132	=>	145,
		50133	=>	145,
		50134	=>	145,
		50135	=>	145,
		50136	=>	146,
		50137	=>	146,
		50138	=>	146,
		50139	=>	147,
		50140	=>	147,
		50141	=>	147,
		50142	=>	147,
		50143	=>	148,
		50144	=>	148,
		50145	=>	148,
		50146	=>	149,
		50147	=>	149,
		50148	=>	149,
		50149	=>	150,
		50150	=>	150,
		50151	=>	150,
		50152	=>	150,
		50153	=>	151,
		50154	=>	151,
		50155	=>	151,
		50156	=>	152,
		50157	=>	152,
		50158	=>	152,
		50159	=>	153,
		50160	=>	153,
		50161	=>	153,
		50162	=>	154,
		50163	=>	154,
		50164	=>	154,
		50165	=>	154,
		50166	=>	155,
		50167	=>	155,
		50168	=>	155,
		50169	=>	156,
		50170	=>	156,
		50171	=>	156,
		50172	=>	157,
		50173	=>	157,
		50174	=>	157,
		50175	=>	157,
		50176	=>	158,
		50177	=>	158,
		50178	=>	158,
		50179	=>	159,
		50180	=>	159,
		50181	=>	159,
		50182	=>	160,
		50183	=>	160,
		50184	=>	160,
		50185	=>	161,
		50186	=>	161,
		50187	=>	161,
		50188	=>	162,
		50189	=>	162,
		50190	=>	162,
		50191	=>	162,
		50192	=>	163,
		50193	=>	163,
		50194	=>	163,
		50195	=>	164,
		50196	=>	164,
		50197	=>	164,
		50198	=>	165,
		50199	=>	165,
		50200	=>	165,
		50201	=>	166,
		50202	=>	166,
		50203	=>	166,
		50204	=>	167,
		50205	=>	167,
		50206	=>	167,
		50207	=>	167,
		50208	=>	168,
		50209	=>	168,
		50210	=>	168,
		50211	=>	169,
		50212	=>	169,
		50213	=>	169,
		50214	=>	170,
		50215	=>	170,
		50216	=>	170,
		50217	=>	171,
		50218	=>	171,
		50219	=>	171,
		50220	=>	172,
		50221	=>	172,
		50222	=>	172,
		50223	=>	173,
		50224	=>	173,
		50225	=>	173,
		50226	=>	174,
		50227	=>	174,
		50228	=>	174,
		50229	=>	175,
		50230	=>	175,
		50231	=>	175,
		50232	=>	175,
		50233	=>	176,
		50234	=>	176,
		50235	=>	176,
		50236	=>	177,
		50237	=>	177,
		50238	=>	177,
		50239	=>	178,
		50240	=>	178,
		50241	=>	178,
		50242	=>	179,
		50243	=>	179,
		50244	=>	179,
		50245	=>	180,
		50246	=>	180,
		50247	=>	180,
		50248	=>	181,
		50249	=>	181,
		50250	=>	181,
		50251	=>	182,
		50252	=>	182,
		50253	=>	182,
		50254	=>	183,
		50255	=>	183,
		50256	=>	183,
		50257	=>	184,
		50258	=>	184,
		50259	=>	184,
		50260	=>	185,
		50261	=>	185,
		50262	=>	185,
		50263	=>	186,
		50264	=>	186,
		50265	=>	186,
		50266	=>	187,
		50267	=>	187,
		50268	=>	187,
		50269	=>	188,
		50270	=>	188,
		50271	=>	188,
		50272	=>	189,
		50273	=>	189,
		50274	=>	189,
		50275	=>	190,
		50276	=>	190,
		50277	=>	190,
		50278	=>	191,
		50279	=>	191,
		50280	=>	191,
		50281	=>	192,
		50282	=>	192,
		50283	=>	192,
		50284	=>	193,
		50285	=>	193,
		50286	=>	193,
		50287	=>	194,
		50288	=>	194,
		50289	=>	194,
		50290	=>	195,
		50291	=>	195,
		50292	=>	196,
		50293	=>	196,
		50294	=>	196,
		50295	=>	197,
		50296	=>	197,
		50297	=>	197,
		50298	=>	198,
		50299	=>	198,
		50300	=>	198,
		50301	=>	199,
		50302	=>	199,
		50303	=>	199,
		50304	=>	200,
		50305	=>	200,
		50306	=>	200,
		50307	=>	201,
		50308	=>	201,
		50309	=>	201,
		50310	=>	202,
		50311	=>	202,
		50312	=>	202,
		50313	=>	203,
		50314	=>	203,
		50315	=>	203,
		50316	=>	204,
		50317	=>	204,
		50318	=>	205,
		50319	=>	205,
		50320	=>	205,
		50321	=>	206,
		50322	=>	206,
		50323	=>	206,
		50324	=>	207,
		50325	=>	207,
		50326	=>	207,
		50327	=>	208,
		50328	=>	208,
		50329	=>	208,
		50330	=>	209,
		50331	=>	209,
		50332	=>	209,
		50333	=>	210,
		50334	=>	210,
		50335	=>	211,
		50336	=>	211,
		50337	=>	211,
		50338	=>	212,
		50339	=>	212,
		50340	=>	212,
		50341	=>	213,
		50342	=>	213,
		50343	=>	213,
		50344	=>	214,
		50345	=>	214,
		50346	=>	214,
		50347	=>	215,
		50348	=>	215,
		50349	=>	216,
		50350	=>	216,
		50351	=>	216,
		50352	=>	217,
		50353	=>	217,
		50354	=>	217,
		50355	=>	218,
		50356	=>	218,
		50357	=>	218,
		50358	=>	219,
		50359	=>	219,
		50360	=>	220,
		50361	=>	220,
		50362	=>	220,
		50363	=>	221,
		50364	=>	221,
		50365	=>	221,
		50366	=>	222,
		50367	=>	222,
		50368	=>	222,
		50369	=>	223,
		50370	=>	223,
		50371	=>	224,
		50372	=>	224,
		50373	=>	224,
		50374	=>	225,
		50375	=>	225,
		50376	=>	225,
		50377	=>	226,
		50378	=>	226,
		50379	=>	226,
		50380	=>	227,
		50381	=>	227,
		50382	=>	228,
		50383	=>	228,
		50384	=>	228,
		50385	=>	229,
		50386	=>	229,
		50387	=>	229,
		50388	=>	230,
		50389	=>	230,
		50390	=>	231,
		50391	=>	231,
		50392	=>	231,
		50393	=>	232,
		50394	=>	232,
		50395	=>	232,
		50396	=>	233,
		50397	=>	233,
		50398	=>	234,
		50399	=>	234,
		50400	=>	234,
		50401	=>	235,
		50402	=>	235,
		50403	=>	235,
		50404	=>	236,
		50405	=>	236,
		50406	=>	237,
		50407	=>	237,
		50408	=>	237,
		50409	=>	238,
		50410	=>	238,
		50411	=>	238,
		50412	=>	239,
		50413	=>	239,
		50414	=>	240,
		50415	=>	240,
		50416	=>	240,
		50417	=>	241,
		50418	=>	241,
		50419	=>	241,
		50420	=>	242,
		50421	=>	242,
		50422	=>	243,
		50423	=>	243,
		50424	=>	243,
		50425	=>	244,
		50426	=>	244,
		50427	=>	245,
		50428	=>	245,
		50429	=>	245,
		50430	=>	246,
		50431	=>	246,
		50432	=>	246,
		50433	=>	247,
		50434	=>	247,
		50435	=>	248,
		50436	=>	248,
		50437	=>	248,
		50438	=>	249,
		50439	=>	249,
		50440	=>	250,
		50441	=>	250,
		50442	=>	250,
		50443	=>	251,
		50444	=>	251,
		50445	=>	251,
		50446	=>	252,
		50447	=>	252,
		50448	=>	253,
		50449	=>	253,
		50450	=>	253,
		50451	=>	254,
		50452	=>	254,
		50453	=>	255,
		50454	=>	255,
		50455	=>	255,
		50456	=>	256,
		50457	=>	256,
		50458	=>	257,
		50459	=>	257,
		50460	=>	257,
		50461	=>	258,
		50462	=>	258,
		50463	=>	258,
		50464	=>	259,
		50465	=>	259,
		50466	=>	260,
		50467	=>	260,
		50468	=>	260,
		50469	=>	261,
		50470	=>	261,
		50471	=>	262,
		50472	=>	262,
		50473	=>	262,
		50474	=>	263,
		50475	=>	263,
		50476	=>	264,
		50477	=>	264,
		50478	=>	264,
		50479	=>	265,
		50480	=>	265,
		50481	=>	266,
		50482	=>	266,
		50483	=>	266,
		50484	=>	267,
		50485	=>	267,
		50486	=>	268,
		50487	=>	268,
		50488	=>	268,
		50489	=>	269,
		50490	=>	269,
		50491	=>	270,
		50492	=>	270,
		50493	=>	270,
		50494	=>	271,
		50495	=>	271,
		50496	=>	272,
		50497	=>	272,
		50498	=>	272,
		50499	=>	273,
		50500	=>	273,
		50501	=>	274,
		50502	=>	274,
		50503	=>	274,
		50504	=>	275,
		50505	=>	275,
		50506	=>	276,
		50507	=>	276,
		50508	=>	277,
		50509	=>	277,
		50510	=>	277,
		50511	=>	278,
		50512	=>	278,
		50513	=>	279,
		50514	=>	279,
		50515	=>	279,
		50516	=>	280,
		50517	=>	280,
		50518	=>	281,
		50519	=>	281,
		50520	=>	281,
		50521	=>	282,
		50522	=>	282,
		50523	=>	283,
		50524	=>	283,
		50525	=>	283,
		50526	=>	284,
		50527	=>	284,
		50528	=>	285,
		50529	=>	285,
		50530	=>	286,
		50531	=>	286,
		50532	=>	286,
		50533	=>	287,
		50534	=>	287,
		50535	=>	288,
		50536	=>	288,
		50537	=>	288,
		50538	=>	289,
		50539	=>	289,
		50540	=>	290,
		50541	=>	290,
		50542	=>	291,
		50543	=>	291,
		50544	=>	291,
		50545	=>	292,
		50546	=>	292,
		50547	=>	293,
		50548	=>	293,
		50549	=>	293,
		50550	=>	294,
		50551	=>	294,
		50552	=>	295,
		50553	=>	295,
		50554	=>	296,
		50555	=>	296,
		50556	=>	296,
		50557	=>	297,
		50558	=>	297,
		50559	=>	298,
		50560	=>	298,
		50561	=>	299,
		50562	=>	299,
		50563	=>	299,
		50564	=>	300,
		50565	=>	300,
		50566	=>	301,
		50567	=>	301,
		50568	=>	301,
		50569	=>	302,
		50570	=>	302,
		50571	=>	303,
		50572	=>	303,
		50573	=>	304,
		50574	=>	304,
		50575	=>	304,
		50576	=>	305,
		50577	=>	305,
		50578	=>	306,
		50579	=>	306,
		50580	=>	307,
		50581	=>	307,
		50582	=>	307,
		50583	=>	308,
		50584	=>	308,
		50585	=>	309,
		50586	=>	309,
		50587	=>	310,
		50588	=>	310,
		50589	=>	310,
		50590	=>	311,
		50591	=>	311,
		50592	=>	312,
		50593	=>	312,
		50594	=>	313,
		50595	=>	313,
		50596	=>	314,
		50597	=>	314,
		50598	=>	314,
		50599	=>	315,
		50600	=>	315,
		50601	=>	316,
		50602	=>	316,
		50603	=>	317,
		50604	=>	317,
		50605	=>	317,
		50606	=>	318,
		50607	=>	318,
		50608	=>	319,
		50609	=>	319,
		50610	=>	320,
		50611	=>	320,
		50612	=>	320,
		50613	=>	321,
		50614	=>	321,
		50615	=>	322,
		50616	=>	322,
		50617	=>	323,
		50618	=>	323,
		50619	=>	324,
		50620	=>	324,
		50621	=>	324,
		50622	=>	325,
		50623	=>	325,
		50624	=>	326,
		50625	=>	326,
		50626	=>	327,
		50627	=>	327,
		50628	=>	328,
		50629	=>	328,
		50630	=>	328,
		50631	=>	329,
		50632	=>	329,
		50633	=>	330,
		50634	=>	330,
		50635	=>	331,
		50636	=>	331,
		50637	=>	332,
		50638	=>	332,
		50639	=>	332,
		50640	=>	333,
		50641	=>	333,
		50642	=>	334,
		50643	=>	334,
		50644	=>	335,
		50645	=>	335,
		50646	=>	336,
		50647	=>	336,
		50648	=>	336,
		50649	=>	337,
		50650	=>	337,
		50651	=>	338,
		50652	=>	338,
		50653	=>	339,
		50654	=>	339,
		50655	=>	340,
		50656	=>	340,
		50657	=>	341,
		50658	=>	341,
		50659	=>	341,
		50660	=>	342,
		50661	=>	342,
		50662	=>	343,
		50663	=>	343,
		50664	=>	344,
		50665	=>	344,
		50666	=>	345,
		50667	=>	345,
		50668	=>	345,
		50669	=>	346,
		50670	=>	346,
		50671	=>	347,
		50672	=>	347,
		50673	=>	348,
		50674	=>	348,
		50675	=>	349,
		50676	=>	349,
		50677	=>	350,
		50678	=>	350,
		50679	=>	351,
		50680	=>	351,
		50681	=>	351,
		50682	=>	352,
		50683	=>	352,
		50684	=>	353,
		50685	=>	353,
		50686	=>	354,
		50687	=>	354,
		50688	=>	355,
		50689	=>	355,
		50690	=>	356,
		50691	=>	356,
		50692	=>	357,
		50693	=>	357,
		50694	=>	357,
		50695	=>	358,
		50696	=>	358,
		50697	=>	359,
		50698	=>	359,
		50699	=>	360,
		50700	=>	360,
		50701	=>	361,
		50702	=>	361,
		50703	=>	362,
		50704	=>	362,
		50705	=>	363,
		50706	=>	363,
		50707	=>	363,
		50708	=>	364,
		50709	=>	364,
		50710	=>	365,
		50711	=>	365,
		50712	=>	366,
		50713	=>	366,
		50714	=>	367,
		50715	=>	367,
		50716	=>	368,
		50717	=>	368,
		50718	=>	369,
		50719	=>	369,
		50720	=>	370,
		50721	=>	370,
		50722	=>	371,
		50723	=>	371,
		50724	=>	371,
		50725	=>	372,
		50726	=>	372,
		50727	=>	373,
		50728	=>	373,
		50729	=>	374,
		50730	=>	374,
		50731	=>	375,
		50732	=>	375,
		50733	=>	376,
		50734	=>	376,
		50735	=>	377,
		50736	=>	377,
		50737	=>	378,
		50738	=>	378,
		50739	=>	379,
		50740	=>	379,
		50741	=>	380,
		50742	=>	380,
		50743	=>	380,
		50744	=>	381,
		50745	=>	381,
		50746	=>	382,
		50747	=>	382,
		50748	=>	383,
		50749	=>	383,
		50750	=>	384,
		50751	=>	384,
		50752	=>	385,
		50753	=>	385,
		50754	=>	386,
		50755	=>	386,
		50756	=>	387,
		50757	=>	387,
		50758	=>	388,
		50759	=>	388,
		50760	=>	389,
		50761	=>	389,
		50762	=>	390,
		50763	=>	390,
		50764	=>	391,
		50765	=>	391,
		50766	=>	392,
		50767	=>	392,
		50768	=>	392,
		50769	=>	393,
		50770	=>	393,
		50771	=>	394,
		50772	=>	394,
		50773	=>	395,
		50774	=>	395,
		50775	=>	396,
		50776	=>	396,
		50777	=>	397,
		50778	=>	397,
		50779	=>	398,
		50780	=>	398,
		50781	=>	399,
		50782	=>	399,
		50783	=>	400,
		50784	=>	400,
		50785	=>	401,
		50786	=>	401,
		50787	=>	402,
		50788	=>	402,
		50789	=>	403,
		50790	=>	403,
		50791	=>	404,
		50792	=>	404,
		50793	=>	405,
		50794	=>	405,
		50795	=>	406,
		50796	=>	406,
		50797	=>	407,
		50798	=>	407,
		50799	=>	408,
		50800	=>	408,
		50801	=>	409,
		50802	=>	409,
		50803	=>	410,
		50804	=>	410,
		50805	=>	411,
		50806	=>	411,
		50807	=>	412,
		50808	=>	412,
		50809	=>	413,
		50810	=>	413,
		50811	=>	414,
		50812	=>	414,
		50813	=>	415,
		50814	=>	415,
		50815	=>	416,
		50816	=>	416,
		50817	=>	417,
		50818	=>	417,
		50819	=>	418,
		50820	=>	418,
		50821	=>	419,
		50822	=>	419,
		50823	=>	420,
		50824	=>	420,
		50825	=>	421,
		50826	=>	421,
		50827	=>	422,
		50828	=>	422,
		50829	=>	423,
		50830	=>	423,
		50831	=>	424,
		50832	=>	424,
		50833	=>	425,
		50834	=>	425,
		50835	=>	426,
		50836	=>	426,
		50837	=>	427,
		50838	=>	427,
		50839	=>	428,
		50840	=>	428,
		50841	=>	429,
		50842	=>	429,
		50843	=>	430,
		50844	=>	430,
		50845	=>	431,
		50846	=>	431,
		50847	=>	432,
		50848	=>	432,
		50849	=>	433,
		50850	=>	433,
		50851	=>	434,
		50852	=>	434,
		50853	=>	435,
		50854	=>	435,
		50855	=>	436,
		50856	=>	436,
		50857	=>	437,
		50858	=>	437,
		50859	=>	438,
		50860	=>	438,
		50861	=>	439,
		50862	=>	439,
		50863	=>	440,
		50864	=>	440,
		50865	=>	441,
		50866	=>	441,
		50867	=>	442,
		50868	=>	442,
		50869	=>	443,
		50870	=>	443,
		50871	=>	444,
		50872	=>	445,
		50873	=>	445,
		50874	=>	446,
		50875	=>	446,
		50876	=>	447,
		50877	=>	447,
		50878	=>	448,
		50879	=>	448,
		50880	=>	449,
		50881	=>	449,
		50882	=>	450,
		50883	=>	450,
		50884	=>	451,
		50885	=>	451,
		50886	=>	452,
		50887	=>	452,
		50888	=>	453,
		50889	=>	453,
		50890	=>	454,
		50891	=>	454,
		50892	=>	455,
		50893	=>	455,
		50894	=>	456,
		50895	=>	456,
		50896	=>	457,
		50897	=>	457,
		50898	=>	458,
		50899	=>	459,
		50900	=>	459,
		50901	=>	460,
		50902	=>	460,
		50903	=>	461,
		50904	=>	461,
		50905	=>	462,
		50906	=>	462,
		50907	=>	463,
		50908	=>	463,
		50909	=>	464,
		50910	=>	464,
		50911	=>	465,
		50912	=>	465,
		50913	=>	466,
		50914	=>	466,
		50915	=>	467,
		50916	=>	467,
		50917	=>	468,
		50918	=>	469,
		50919	=>	469,
		50920	=>	470,
		50921	=>	470,
		50922	=>	471,
		50923	=>	471,
		50924	=>	472,
		50925	=>	472,
		50926	=>	473,
		50927	=>	473,
		50928	=>	474,
		50929	=>	474,
		50930	=>	475,
		50931	=>	475,
		50932	=>	476,
		50933	=>	477,
		50934	=>	477,
		50935	=>	478,
		50936	=>	478,
		50937	=>	479,
		50938	=>	479,
		50939	=>	480,
		50940	=>	480,
		50941	=>	481,
		50942	=>	481,
		50943	=>	482,
		50944	=>	482,
		50945	=>	483,
		50946	=>	483,
		50947	=>	484,
		50948	=>	485,
		50949	=>	485,
		50950	=>	486,
		50951	=>	486,
		50952	=>	487,
		50953	=>	487,
		50954	=>	488,
		50955	=>	488,
		50956	=>	489,
		50957	=>	489,
		50958	=>	490,
		50959	=>	491,
		50960	=>	491,
		50961	=>	492,
		50962	=>	492,
		50963	=>	493,
		50964	=>	493,
		50965	=>	494,
		50966	=>	494,
		50967	=>	495,
		50968	=>	495,
		50969	=>	496,
		50970	=>	496,
		50971	=>	497,
		50972	=>	498,
		50973	=>	498,
		50974	=>	499,
		50975	=>	499,
		50976	=>	500,
		50977	=>	500,
		50978	=>	501,
		50979	=>	501,
		50980	=>	502,
		50981	=>	502,
		50982	=>	503,
		50983	=>	504,
		50984	=>	504,
		50985	=>	505,
		50986	=>	505,
		50987	=>	506,
		50988	=>	506,
		50989	=>	507,
		50990	=>	507,
		50991	=>	508,
		50992	=>	509,
		50993	=>	509,
		50994	=>	510,
		50995	=>	510,
		50996	=>	511,
		50997	=>	511,
		50998	=>	512,
		50999	=>	512,
		51000	=>	513,
		51001	=>	514,
		51002	=>	514,
		51003	=>	515,
		51004	=>	515,
		51005	=>	516,
		51006	=>	516,
		51007	=>	517,
		51008	=>	517,
		51009	=>	518,
		51010	=>	519,
		51011	=>	519,
		51012	=>	520,
		51013	=>	520,
		51014	=>	521,
		51015	=>	521,
		51016	=>	522,
		51017	=>	522,
		51018	=>	523,
		51019	=>	524,
		51020	=>	524,
		51021	=>	525,
		51022	=>	525,
		51023	=>	526,
		51024	=>	526,
		51025	=>	527,
		51026	=>	527,
		51027	=>	528,
		51028	=>	529,
		51029	=>	529,
		51030	=>	530,
		51031	=>	530,
		51032	=>	531,
		51033	=>	531,
		51034	=>	532,
		51035	=>	533,
		51036	=>	533,
		51037	=>	534,
		51038	=>	534,
		51039	=>	535,
		51040	=>	535,
		51041	=>	536,
		51042	=>	536,
		51043	=>	537,
		51044	=>	538,
		51045	=>	538,
		51046	=>	539,
		51047	=>	539,
		51048	=>	540,
		51049	=>	540,
		51050	=>	541,
		51051	=>	542,
		51052	=>	542,
		51053	=>	543,
		51054	=>	543,
		51055	=>	544,
		51056	=>	544,
		51057	=>	545,
		51058	=>	546,
		51059	=>	546,
		51060	=>	547,
		51061	=>	547,
		51062	=>	548,
		51063	=>	548,
		51064	=>	549,
		51065	=>	550,
		51066	=>	550,
		51067	=>	551,
		51068	=>	551,
		51069	=>	552,
		51070	=>	552,
		51071	=>	553,
		51072	=>	554,
		51073	=>	554,
		51074	=>	555,
		51075	=>	555,
		51076	=>	556,
		51077	=>	556,
		51078	=>	557,
		51079	=>	558,
		51080	=>	558,
		51081	=>	559,
		51082	=>	559,
		51083	=>	560,
		51084	=>	561,
		51085	=>	561,
		51086	=>	562,
		51087	=>	562,
		51088	=>	563,
		51089	=>	563,
		51090	=>	564,
		51091	=>	565,
		51092	=>	565,
		51093	=>	566,
		51094	=>	566,
		51095	=>	567,
		51096	=>	567,
		51097	=>	568,
		51098	=>	569,
		51099	=>	569,
		51100	=>	570,
		51101	=>	570,
		51102	=>	571,
		51103	=>	572,
		51104	=>	572,
		51105	=>	573,
		51106	=>	573,
		51107	=>	574,
		51108	=>	574,
		51109	=>	575,
		51110	=>	576,
		51111	=>	576,
		51112	=>	577,
		51113	=>	577,
		51114	=>	578,
		51115	=>	579,
		51116	=>	579,
		51117	=>	580,
		51118	=>	580,
		51119	=>	581,
		51120	=>	582,
		51121	=>	582,
		51122	=>	583,
		51123	=>	583,
		51124	=>	584,
		51125	=>	584,
		51126	=>	585,
		51127	=>	586,
		51128	=>	586,
		51129	=>	587,
		51130	=>	587,
		51131	=>	588,
		51132	=>	589,
		51133	=>	589,
		51134	=>	590,
		51135	=>	590,
		51136	=>	591,
		51137	=>	592,
		51138	=>	592,
		51139	=>	593,
		51140	=>	593,
		51141	=>	594,
		51142	=>	595,
		51143	=>	595,
		51144	=>	596,
		51145	=>	596,
		51146	=>	597,
		51147	=>	598,
		51148	=>	598,
		51149	=>	599,
		51150	=>	599,
		51151	=>	600,
		51152	=>	601,
		51153	=>	601,
		51154	=>	602,
		51155	=>	602,
		51156	=>	603,
		51157	=>	604,
		51158	=>	604,
		51159	=>	605,
		51160	=>	605,
		51161	=>	606,
		51162	=>	607,
		51163	=>	607,
		51164	=>	608,
		51165	=>	608,
		51166	=>	609,
		51167	=>	610,
		51168	=>	610,
		51169	=>	611,
		51170	=>	611,
		51171	=>	612,
		51172	=>	613,
		51173	=>	613,
		51174	=>	614,
		51175	=>	614,
		51176	=>	615,
		51177	=>	616,
		51178	=>	616,
		51179	=>	617,
		51180	=>	617,
		51181	=>	618,
		51182	=>	619,
		51183	=>	619,
		51184	=>	620,
		51185	=>	620,
		51186	=>	621,
		51187	=>	622,
		51188	=>	622,
		51189	=>	623,
		51190	=>	624,
		51191	=>	624,
		51192	=>	625,
		51193	=>	625,
		51194	=>	626,
		51195	=>	627,
		51196	=>	627,
		51197	=>	628,
		51198	=>	628,
		51199	=>	629,
		51200	=>	630,
		51201	=>	630,
		51202	=>	631,
		51203	=>	631,
		51204	=>	632,
		51205	=>	633,
		51206	=>	633,
		51207	=>	634,
		51208	=>	635,
		51209	=>	635,
		51210	=>	636,
		51211	=>	636,
		51212	=>	637,
		51213	=>	638,
		51214	=>	638,
		51215	=>	639,
		51216	=>	639,
		51217	=>	640,
		51218	=>	641,
		51219	=>	641,
		51220	=>	642,
		51221	=>	643,
		51222	=>	643,
		51223	=>	644,
		51224	=>	644,
		51225	=>	645,
		51226	=>	646,
		51227	=>	646,
		51228	=>	647,
		51229	=>	648,
		51230	=>	648,
		51231	=>	649,
		51232	=>	649,
		51233	=>	650,
		51234	=>	651,
		51235	=>	651,
		51236	=>	652,
		51237	=>	652,
		51238	=>	653,
		51239	=>	654,
		51240	=>	654,
		51241	=>	655,
		51242	=>	656,
		51243	=>	656,
		51244	=>	657,
		51245	=>	657,
		51246	=>	658,
		51247	=>	659,
		51248	=>	659,
		51249	=>	660,
		51250	=>	661,
		51251	=>	661,
		51252	=>	662,
		51253	=>	663,
		51254	=>	663,
		51255	=>	664,
		51256	=>	664,
		51257	=>	665,
		51258	=>	666,
		51259	=>	666,
		51260	=>	667,
		51261	=>	668,
		51262	=>	668,
		51263	=>	669,
		51264	=>	669,
		51265	=>	670,
		51266	=>	671,
		51267	=>	671,
		51268	=>	672,
		51269	=>	673,
		51270	=>	673,
		51271	=>	674,
		51272	=>	675,
		51273	=>	675,
		51274	=>	676,
		51275	=>	676,
		51276	=>	677,
		51277	=>	678,
		51278	=>	678,
		51279	=>	679,
		51280	=>	680,
		51281	=>	680,
		51282	=>	681,
		51283	=>	682,
		51284	=>	682,
		51285	=>	683,
		51286	=>	683,
		51287	=>	684,
		51288	=>	685,
		51289	=>	685,
		51290	=>	686,
		51291	=>	687,
		51292	=>	687,
		51293	=>	688,
		51294	=>	689,
		51295	=>	689,
		51296	=>	690,
		51297	=>	690,
		51298	=>	691,
		51299	=>	692,
		51300	=>	692,
		51301	=>	693,
		51302	=>	694,
		51303	=>	694,
		51304	=>	695,
		51305	=>	696,
		51306	=>	696,
		51307	=>	697,
		51308	=>	698,
		51309	=>	698,
		51310	=>	699,
		51311	=>	699,
		51312	=>	700,
		51313	=>	701,
		51314	=>	701,
		51315	=>	702,
		51316	=>	703,
		51317	=>	703,
		51318	=>	704,
		51319	=>	705,
		51320	=>	705,
		51321	=>	706,
		51322	=>	707,
		51323	=>	707,
		51324	=>	708,
		51325	=>	709,
		51326	=>	709,
		51327	=>	710,
		51328	=>	710,
		51329	=>	711,
		51330	=>	712,
		51331	=>	712,
		51332	=>	713,
		51333	=>	714,
		51334	=>	714,
		51335	=>	715,
		51336	=>	716,
		51337	=>	716,
		51338	=>	717,
		51339	=>	718,
		51340	=>	718,
		51341	=>	719,
		51342	=>	720,
		51343	=>	720,
		51344	=>	721,
		51345	=>	722,
		51346	=>	722,
		51347	=>	723,
		51348	=>	724,
		51349	=>	724,
		51350	=>	725,
		51351	=>	726,
		51352	=>	726,
		51353	=>	727,
		51354	=>	728,
		51355	=>	728,
		51356	=>	729,
		51357	=>	729,
		51358	=>	730,
		51359	=>	731,
		51360	=>	731,
		51361	=>	732,
		51362	=>	733,
		51363	=>	733,
		51364	=>	734,
		51365	=>	735,
		51366	=>	735,
		51367	=>	736,
		51368	=>	737,
		51369	=>	737,
		51370	=>	738,
		51371	=>	739,
		51372	=>	739,
		51373	=>	740,
		51374	=>	741,
		51375	=>	741,
		51376	=>	742,
		51377	=>	743,
		51378	=>	743,
		51379	=>	744,
		51380	=>	745,
		51381	=>	745,
		51382	=>	746,
		51383	=>	747,
		51384	=>	747,
		51385	=>	748,
		51386	=>	749,
		51387	=>	749,
		51388	=>	750,
		51389	=>	751,
		51390	=>	751,
		51391	=>	752,
		51392	=>	753,
		51393	=>	753,
		51394	=>	754,
		51395	=>	755,
		51396	=>	755,
		51397	=>	756,
		51398	=>	757,
		51399	=>	757,
		51400	=>	758,
		51401	=>	759,
		51402	=>	759,
		51403	=>	760,
		51404	=>	761,
		51405	=>	761,
		51406	=>	762,
		51407	=>	763,
		51408	=>	763,
		51409	=>	764,
		51410	=>	765,
		51411	=>	766,
		51412	=>	766,
		51413	=>	767,
		51414	=>	768,
		51415	=>	768,
		51416	=>	769,
		51417	=>	770,
		51418	=>	770,
		51419	=>	771,
		51420	=>	772,
		51421	=>	772,
		51422	=>	773,
		51423	=>	774,
		51424	=>	774,
		51425	=>	775,
		51426	=>	776,
		51427	=>	776,
		51428	=>	777,
		51429	=>	778,
		51430	=>	778,
		51431	=>	779,
		51432	=>	780,
		51433	=>	780,
		51434	=>	781,
		51435	=>	782,
		51436	=>	782,
		51437	=>	783,
		51438	=>	784,
		51439	=>	785,
		51440	=>	785,
		51441	=>	786,
		51442	=>	787,
		51443	=>	787,
		51444	=>	788,
		51445	=>	789,
		51446	=>	789,
		51447	=>	790,
		51448	=>	791,
		51449	=>	791,
		51450	=>	792,
		51451	=>	793,
		51452	=>	793,
		51453	=>	794,
		51454	=>	795,
		51455	=>	795,
		51456	=>	796,
		51457	=>	797,
		51458	=>	798,
		51459	=>	798,
		51460	=>	799,
		51461	=>	800,
		51462	=>	800,
		51463	=>	801,
		51464	=>	802,
		51465	=>	802,
		51466	=>	803,
		51467	=>	804,
		51468	=>	804,
		51469	=>	805,
		51470	=>	806,
		51471	=>	807,
		51472	=>	807,
		51473	=>	808,
		51474	=>	809,
		51475	=>	809,
		51476	=>	810,
		51477	=>	811,
		51478	=>	811,
		51479	=>	812,
		51480	=>	813,
		51481	=>	813,
		51482	=>	814,
		51483	=>	815,
		51484	=>	816,
		51485	=>	816,
		51486	=>	817,
		51487	=>	818,
		51488	=>	818,
		51489	=>	819,
		51490	=>	820,
		51491	=>	820,
		51492	=>	821,
		51493	=>	822,
		51494	=>	823,
		51495	=>	823,
		51496	=>	824,
		51497	=>	825,
		51498	=>	825,
		51499	=>	826,
		51500	=>	827,
		51501	=>	827,
		51502	=>	828,
		51503	=>	829,
		51504	=>	830,
		51505	=>	830,
		51506	=>	831,
		51507	=>	832,
		51508	=>	832,
		51509	=>	833,
		51510	=>	834,
		51511	=>	834,
		51512	=>	835,
		51513	=>	836,
		51514	=>	837,
		51515	=>	837,
		51516	=>	838,
		51517	=>	839,
		51518	=>	839,
		51519	=>	840,
		51520	=>	841,
		51521	=>	842,
		51522	=>	842,
		51523	=>	843,
		51524	=>	844,
		51525	=>	844,
		51526	=>	845,
		51527	=>	846,
		51528	=>	847,
		51529	=>	847,
		51530	=>	848,
		51531	=>	849,
		51532	=>	849,
		51533	=>	850,
		51534	=>	851,
		51535	=>	851,
		51536	=>	852,
		51537	=>	853,
		51538	=>	854,
		51539	=>	854,
		51540	=>	855,
		51541	=>	856,
		51542	=>	856,
		51543	=>	857,
		51544	=>	858,
		51545	=>	859,
		51546	=>	859,
		51547	=>	860,
		51548	=>	861,
		51549	=>	861,
		51550	=>	862,
		51551	=>	863,
		51552	=>	864,
		51553	=>	864,
		51554	=>	865,
		51555	=>	866,
		51556	=>	866,
		51557	=>	867,
		51558	=>	868,
		51559	=>	869,
		51560	=>	869,
		51561	=>	870,
		51562	=>	871,
		51563	=>	872,
		51564	=>	872,
		51565	=>	873,
		51566	=>	874,
		51567	=>	874,
		51568	=>	875,
		51569	=>	876,
		51570	=>	877,
		51571	=>	877,
		51572	=>	878,
		51573	=>	879,
		51574	=>	879,
		51575	=>	880,
		51576	=>	881,
		51577	=>	882,
		51578	=>	882,
		51579	=>	883,
		51580	=>	884,
		51581	=>	885,
		51582	=>	885,
		51583	=>	886,
		51584	=>	887,
		51585	=>	887,
		51586	=>	888,
		51587	=>	889,
		51588	=>	890,
		51589	=>	890,
		51590	=>	891,
		51591	=>	892,
		51592	=>	893,
		51593	=>	893,
		51594	=>	894,
		51595	=>	895,
		51596	=>	895,
		51597	=>	896,
		51598	=>	897,
		51599	=>	898,
		51600	=>	898,
		51601	=>	899,
		51602	=>	900,
		51603	=>	901,
		51604	=>	901,
		51605	=>	902,
		51606	=>	903,
		51607	=>	903,
		51608	=>	904,
		51609	=>	905,
		51610	=>	906,
		51611	=>	906,
		51612	=>	907,
		51613	=>	908,
		51614	=>	909,
		51615	=>	909,
		51616	=>	910,
		51617	=>	911,
		51618	=>	912,
		51619	=>	912,
		51620	=>	913,
		51621	=>	914,
		51622	=>	914,
		51623	=>	915,
		51624	=>	916,
		51625	=>	917,
		51626	=>	917,
		51627	=>	918,
		51628	=>	919,
		51629	=>	920,
		51630	=>	920,
		51631	=>	921,
		51632	=>	922,
		51633	=>	923,
		51634	=>	923,
		51635	=>	924,
		51636	=>	925,
		51637	=>	926,
		51638	=>	926,
		51639	=>	927,
		51640	=>	928,
		51641	=>	929,
		51642	=>	929,
		51643	=>	930,
		51644	=>	931,
		51645	=>	932,
		51646	=>	932,
		51647	=>	933,
		51648	=>	934,
		51649	=>	934,
		51650	=>	935,
		51651	=>	936,
		51652	=>	937,
		51653	=>	937,
		51654	=>	938,
		51655	=>	939,
		51656	=>	940,
		51657	=>	940,
		51658	=>	941,
		51659	=>	942,
		51660	=>	943,
		51661	=>	943,
		51662	=>	944,
		51663	=>	945,
		51664	=>	946,
		51665	=>	946,
		51666	=>	947,
		51667	=>	948,
		51668	=>	949,
		51669	=>	949,
		51670	=>	950,
		51671	=>	951,
		51672	=>	952,
		51673	=>	952,
		51674	=>	953,
		51675	=>	954,
		51676	=>	955,
		51677	=>	955,
		51678	=>	956,
		51679	=>	957,
		51680	=>	958,
		51681	=>	958,
		51682	=>	959,
		51683	=>	960,
		51684	=>	961,
		51685	=>	961,
		51686	=>	962,
		51687	=>	963,
		51688	=>	964,
		51689	=>	965,
		51690	=>	965,
		51691	=>	966,
		51692	=>	967,
		51693	=>	968,
		51694	=>	968,
		51695	=>	969,
		51696	=>	970,
		51697	=>	971,
		51698	=>	971,
		51699	=>	972,
		51700	=>	973,
		51701	=>	974,
		51702	=>	974,
		51703	=>	975,
		51704	=>	976,
		51705	=>	977,
		51706	=>	977,
		51707	=>	978,
		51708	=>	979,
		51709	=>	980,
		51710	=>	980,
		51711	=>	981,
		51712	=>	982,
		51713	=>	983,
		51714	=>	984,
		51715	=>	984,
		51716	=>	985,
		51717	=>	986,
		51718	=>	987,
		51719	=>	987,
		51720	=>	988,
		51721	=>	989,
		51722	=>	990,
		51723	=>	990,
		51724	=>	991,
		51725	=>	992,
		51726	=>	993,
		51727	=>	993,
		51728	=>	994,
		51729	=>	995,
		51730	=>	996,
		51731	=>	997,
		51732	=>	997,
		51733	=>	998,
		51734	=>	999,
		51735	=>	1000,
		51736	=>	1000,
		51737	=>	1001,
		51738	=>	1002,
		51739	=>	1003,
		51740	=>	1003,
		51741	=>	1004,
		51742	=>	1005,
		51743	=>	1006,
		51744	=>	1007,
		51745	=>	1007,
		51746	=>	1008,
		51747	=>	1009,
		51748	=>	1010,
		51749	=>	1010,
		51750	=>	1011,
		51751	=>	1012,
		51752	=>	1013,
		51753	=>	1014,
		51754	=>	1014,
		51755	=>	1015,
		51756	=>	1016,
		51757	=>	1017,
		51758	=>	1017,
		51759	=>	1018,
		51760	=>	1019,
		51761	=>	1020,
		51762	=>	1021,
		51763	=>	1021,
		51764	=>	1022,
		51765	=>	1023,
		51766	=>	1024,
		51767	=>	1024,
		51768	=>	1025,
		51769	=>	1026,
		51770	=>	1027,
		51771	=>	1028,
		51772	=>	1028,
		51773	=>	1029,
		51774	=>	1030,
		51775	=>	1031,
		51776	=>	1031,
		51777	=>	1032,
		51778	=>	1033,
		51779	=>	1034,
		51780	=>	1035,
		51781	=>	1035,
		51782	=>	1036,
		51783	=>	1037,
		51784	=>	1038,
		51785	=>	1039,
		51786	=>	1039,
		51787	=>	1040,
		51788	=>	1041,
		51789	=>	1042,
		51790	=>	1042,
		51791	=>	1043,
		51792	=>	1044,
		51793	=>	1045,
		51794	=>	1046,
		51795	=>	1046,
		51796	=>	1047,
		51797	=>	1048,
		51798	=>	1049,
		51799	=>	1050,
		51800	=>	1050,
		51801	=>	1051,
		51802	=>	1052,
		51803	=>	1053,
		51804	=>	1053,
		51805	=>	1054,
		51806	=>	1055,
		51807	=>	1056,
		51808	=>	1057,
		51809	=>	1057,
		51810	=>	1058,
		51811	=>	1059,
		51812	=>	1060,
		51813	=>	1061,
		51814	=>	1061,
		51815	=>	1062,
		51816	=>	1063,
		51817	=>	1064,
		51818	=>	1065,
		51819	=>	1065,
		51820	=>	1066,
		51821	=>	1067,
		51822	=>	1068,
		51823	=>	1069,
		51824	=>	1069,
		51825	=>	1070,
		51826	=>	1071,
		51827	=>	1072,
		51828	=>	1073,
		51829	=>	1073,
		51830	=>	1074,
		51831	=>	1075,
		51832	=>	1076,
		51833	=>	1077,
		51834	=>	1077,
		51835	=>	1078,
		51836	=>	1079,
		51837	=>	1080,
		51838	=>	1080,
		51839	=>	1081,
		51840	=>	1082,
		51841	=>	1083,
		51842	=>	1084,
		51843	=>	1085,
		51844	=>	1085,
		51845	=>	1086,
		51846	=>	1087,
		51847	=>	1088,
		51848	=>	1089,
		51849	=>	1089,
		51850	=>	1090,
		51851	=>	1091,
		51852	=>	1092,
		51853	=>	1093,
		51854	=>	1093,
		51855	=>	1094,
		51856	=>	1095,
		51857	=>	1096,
		51858	=>	1097,
		51859	=>	1097,
		51860	=>	1098,
		51861	=>	1099,
		51862	=>	1100,
		51863	=>	1101,
		51864	=>	1101,
		51865	=>	1102,
		51866	=>	1103,
		51867	=>	1104,
		51868	=>	1105,
		51869	=>	1105,
		51870	=>	1106,
		51871	=>	1107,
		51872	=>	1108,
		51873	=>	1109,
		51874	=>	1109,
		51875	=>	1110,
		51876	=>	1111,
		51877	=>	1112,
		51878	=>	1113,
		51879	=>	1114,
		51880	=>	1114,
		51881	=>	1115,
		51882	=>	1116,
		51883	=>	1117,
		51884	=>	1118,
		51885	=>	1118,
		51886	=>	1119,
		51887	=>	1120,
		51888	=>	1121,
		51889	=>	1122,
		51890	=>	1122,
		51891	=>	1123,
		51892	=>	1124,
		51893	=>	1125,
		51894	=>	1126,
		51895	=>	1127,
		51896	=>	1127,
		51897	=>	1128,
		51898	=>	1129,
		51899	=>	1130,
		51900	=>	1131,
		51901	=>	1131,
		51902	=>	1132,
		51903	=>	1133,
		51904	=>	1134,
		51905	=>	1135,
		51906	=>	1136,
		51907	=>	1136,
		51908	=>	1137,
		51909	=>	1138,
		51910	=>	1139,
		51911	=>	1140,
		51912	=>	1141,
		51913	=>	1141,
		51914	=>	1142,
		51915	=>	1143,
		51916	=>	1144,
		51917	=>	1145,
		51918	=>	1145,
		51919	=>	1146,
		51920	=>	1147,
		51921	=>	1148,
		51922	=>	1149,
		51923	=>	1150,
		51924	=>	1150,
		51925	=>	1151,
		51926	=>	1152,
		51927	=>	1153,
		51928	=>	1154,
		51929	=>	1155,
		51930	=>	1155,
		51931	=>	1156,
		51932	=>	1157,
		51933	=>	1158,
		51934	=>	1159,
		51935	=>	1159,
		51936	=>	1160,
		51937	=>	1161,
		51938	=>	1162,
		51939	=>	1163,
		51940	=>	1164,
		51941	=>	1164,
		51942	=>	1165,
		51943	=>	1166,
		51944	=>	1167,
		51945	=>	1168,
		51946	=>	1169,
		51947	=>	1169,
		51948	=>	1170,
		51949	=>	1171,
		51950	=>	1172,
		51951	=>	1173,
		51952	=>	1174,
		51953	=>	1174,
		51954	=>	1175,
		51955	=>	1176,
		51956	=>	1177,
		51957	=>	1178,
		51958	=>	1179,
		51959	=>	1179,
		51960	=>	1180,
		51961	=>	1181,
		51962	=>	1182,
		51963	=>	1183,
		51964	=>	1184,
		51965	=>	1184,
		51966	=>	1185,
		51967	=>	1186,
		51968	=>	1187,
		51969	=>	1188,
		51970	=>	1189,
		51971	=>	1189,
		51972	=>	1190,
		51973	=>	1191,
		51974	=>	1192,
		51975	=>	1193,
		51976	=>	1194,
		51977	=>	1195,
		51978	=>	1195,
		51979	=>	1196,
		51980	=>	1197,
		51981	=>	1198,
		51982	=>	1199,
		51983	=>	1200,
		51984	=>	1200,
		51985	=>	1201,
		51986	=>	1202,
		51987	=>	1203,
		51988	=>	1204,
		51989	=>	1205,
		51990	=>	1205,
		51991	=>	1206,
		51992	=>	1207,
		51993	=>	1208,
		51994	=>	1209,
		51995	=>	1210,
		51996	=>	1211,
		51997	=>	1211,
		51998	=>	1212,
		51999	=>	1213,
		52000	=>	1214,
		52001	=>	1215,
		52002	=>	1216,
		52003	=>	1216,
		52004	=>	1217,
		52005	=>	1218,
		52006	=>	1219,
		52007	=>	1220,
		52008	=>	1221,
		52009	=>	1222,
		52010	=>	1222,
		52011	=>	1223,
		52012	=>	1224,
		52013	=>	1225,
		52014	=>	1226,
		52015	=>	1227,
		52016	=>	1228,
		52017	=>	1228,
		52018	=>	1229,
		52019	=>	1230,
		52020	=>	1231,
		52021	=>	1232,
		52022	=>	1233,
		52023	=>	1233,
		52024	=>	1234,
		52025	=>	1235,
		52026	=>	1236,
		52027	=>	1237,
		52028	=>	1238,
		52029	=>	1239,
		52030	=>	1239,
		52031	=>	1240,
		52032	=>	1241,
		52033	=>	1242,
		52034	=>	1243,
		52035	=>	1244,
		52036	=>	1245,
		52037	=>	1245,
		52038	=>	1246,
		52039	=>	1247,
		52040	=>	1248,
		52041	=>	1249,
		52042	=>	1250,
		52043	=>	1251,
		52044	=>	1251,
		52045	=>	1252,
		52046	=>	1253,
		52047	=>	1254,
		52048	=>	1255,
		52049	=>	1256,
		52050	=>	1257,
		52051	=>	1258,
		52052	=>	1258,
		52053	=>	1259,
		52054	=>	1260,
		52055	=>	1261,
		52056	=>	1262,
		52057	=>	1263,
		52058	=>	1264,
		52059	=>	1264,
		52060	=>	1265,
		52061	=>	1266,
		52062	=>	1267,
		52063	=>	1268,
		52064	=>	1269,
		52065	=>	1270,
		52066	=>	1270,
		52067	=>	1271,
		52068	=>	1272,
		52069	=>	1273,
		52070	=>	1274,
		52071	=>	1275,
		52072	=>	1276,
		52073	=>	1277,
		52074	=>	1277,
		52075	=>	1278,
		52076	=>	1279,
		52077	=>	1280,
		52078	=>	1281,
		52079	=>	1282,
		52080	=>	1283,
		52081	=>	1284,
		52082	=>	1284,
		52083	=>	1285,
		52084	=>	1286,
		52085	=>	1287,
		52086	=>	1288,
		52087	=>	1289,
		52088	=>	1290,
		52089	=>	1290,
		52090	=>	1291,
		52091	=>	1292,
		52092	=>	1293,
		52093	=>	1294,
		52094	=>	1295,
		52095	=>	1296,
		52096	=>	1297,
		52097	=>	1297,
		52098	=>	1298,
		52099	=>	1299,
		52100	=>	1300,
		52101	=>	1301,
		52102	=>	1302,
		52103	=>	1303,
		52104	=>	1304,
		52105	=>	1304,
		52106	=>	1305,
		52107	=>	1306,
		52108	=>	1307,
		52109	=>	1308,
		52110	=>	1309,
		52111	=>	1310,
		52112	=>	1311,
		52113	=>	1312,
		52114	=>	1312,
		52115	=>	1313,
		52116	=>	1314,
		52117	=>	1315,
		52118	=>	1316,
		52119	=>	1317,
		52120	=>	1318,
		52121	=>	1319,
		52122	=>	1319,
		52123	=>	1320,
		52124	=>	1321,
		52125	=>	1322,
		52126	=>	1323,
		52127	=>	1324,
		52128	=>	1325,
		52129	=>	1326,
		52130	=>	1327,
		52131	=>	1327,
		52132	=>	1328,
		52133	=>	1329,
		52134	=>	1330,
		52135	=>	1331,
		52136	=>	1332,
		52137	=>	1333,
		52138	=>	1334,
		52139	=>	1334,
		52140	=>	1335,
		52141	=>	1336,
		52142	=>	1337,
		52143	=>	1338,
		52144	=>	1339,
		52145	=>	1340,
		52146	=>	1341,
		52147	=>	1342,
		52148	=>	1342,
		52149	=>	1343,
		52150	=>	1344,
		52151	=>	1345,
		52152	=>	1346,
		52153	=>	1347,
		52154	=>	1348,
		52155	=>	1349,
		52156	=>	1350,
		52157	=>	1351,
		52158	=>	1351,
		52159	=>	1352,
		52160	=>	1353,
		52161	=>	1354,
		52162	=>	1355,
		52163	=>	1356,
		52164	=>	1357,
		52165	=>	1358,
		52166	=>	1359,
		52167	=>	1359,
		52168	=>	1360,
		52169	=>	1361,
		52170	=>	1362,
		52171	=>	1363,
		52172	=>	1364,
		52173	=>	1365,
		52174	=>	1366,
		52175	=>	1367,
		52176	=>	1368,
		52177	=>	1368,
		52178	=>	1369,
		52179	=>	1370,
		52180	=>	1371,
		52181	=>	1372,
		52182	=>	1373,
		52183	=>	1374,
		52184	=>	1375,
		52185	=>	1376,
		52186	=>	1377,
		52187	=>	1377,
		52188	=>	1378,
		52189	=>	1379,
		52190	=>	1380,
		52191	=>	1381,
		52192	=>	1382,
		52193	=>	1383,
		52194	=>	1384,
		52195	=>	1385,
		52196	=>	1386,
		52197	=>	1386,
		52198	=>	1387,
		52199	=>	1388,
		52200	=>	1389,
		52201	=>	1390,
		52202	=>	1391,
		52203	=>	1392,
		52204	=>	1393,
		52205	=>	1394,
		52206	=>	1395,
		52207	=>	1395,
		52208	=>	1396,
		52209	=>	1397,
		52210	=>	1398,
		52211	=>	1399,
		52212	=>	1400,
		52213	=>	1401,
		52214	=>	1402,
		52215	=>	1403,
		52216	=>	1404,
		52217	=>	1405,
		52218	=>	1405,
		52219	=>	1406,
		52220	=>	1407,
		52221	=>	1408,
		52222	=>	1409,
		52223	=>	1410,
		52224	=>	1411,
		52225	=>	1412,
		52226	=>	1413,
		52227	=>	1414,
		52228	=>	1415,
		52229	=>	1416,
		52230	=>	1416,
		52231	=>	1417,
		52232	=>	1418,
		52233	=>	1419,
		52234	=>	1420,
		52235	=>	1421,
		52236	=>	1422,
		52237	=>	1423,
		52238	=>	1424,
		52239	=>	1425,
		52240	=>	1426,
		52241	=>	1427,
		52242	=>	1427,
		52243	=>	1428,
		52244	=>	1429,
		52245	=>	1430,
		52246	=>	1431,
		52247	=>	1432,
		52248	=>	1433,
		52249	=>	1434,
		52250	=>	1435,
		52251	=>	1436,
		52252	=>	1437,
		52253	=>	1438,
		52254	=>	1438,
		52255	=>	1439,
		52256	=>	1440,
		52257	=>	1441,
		52258	=>	1442,
		52259	=>	1443,
		52260	=>	1444,
		52261	=>	1445,
		52262	=>	1446,
		52263	=>	1447,
		52264	=>	1448,
		52265	=>	1449,
		52266	=>	1450,
		52267	=>	1450,
		52268	=>	1451,
		52269	=>	1452,
		52270	=>	1453,
		52271	=>	1454,
		52272	=>	1455,
		52273	=>	1456,
		52274	=>	1457,
		52275	=>	1458,
		52276	=>	1459,
		52277	=>	1460,
		52278	=>	1461,
		52279	=>	1462,
		52280	=>	1462,
		52281	=>	1463,
		52282	=>	1464,
		52283	=>	1465,
		52284	=>	1466,
		52285	=>	1467,
		52286	=>	1468,
		52287	=>	1469,
		52288	=>	1470,
		52289	=>	1471,
		52290	=>	1472,
		52291	=>	1473,
		52292	=>	1474,
		52293	=>	1475,
		52294	=>	1475,
		52295	=>	1476,
		52296	=>	1477,
		52297	=>	1478,
		52298	=>	1479,
		52299	=>	1480,
		52300	=>	1481,
		52301	=>	1482,
		52302	=>	1483,
		52303	=>	1484,
		52304	=>	1485,
		52305	=>	1486,
		52306	=>	1487,
		52307	=>	1488,
		52308	=>	1489,
		52309	=>	1490,
		52310	=>	1490,
		52311	=>	1491,
		52312	=>	1492,
		52313	=>	1493,
		52314	=>	1494,
		52315	=>	1495,
		52316	=>	1496,
		52317	=>	1497,
		52318	=>	1498,
		52319	=>	1499,
		52320	=>	1500,
		52321	=>	1501,
		52322	=>	1502,
		52323	=>	1503,
		52324	=>	1504,
		52325	=>	1505,
		52326	=>	1505,
		52327	=>	1506,
		52328	=>	1507,
		52329	=>	1508,
		52330	=>	1509,
		52331	=>	1510,
		52332	=>	1511,
		52333	=>	1512,
		52334	=>	1513,
		52335	=>	1514,
		52336	=>	1515,
		52337	=>	1516,
		52338	=>	1517,
		52339	=>	1518,
		52340	=>	1519,
		52341	=>	1520,
		52342	=>	1521,
		52343	=>	1522,
		52344	=>	1522,
		52345	=>	1523,
		52346	=>	1524,
		52347	=>	1525,
		52348	=>	1526,
		52349	=>	1527,
		52350	=>	1528,
		52351	=>	1529,
		52352	=>	1530,
		52353	=>	1531,
		52354	=>	1532,
		52355	=>	1533,
		52356	=>	1534,
		52357	=>	1535,
		52358	=>	1536,
		52359	=>	1537,
		52360	=>	1538,
		52361	=>	1539,
		52362	=>	1540,
		52363	=>	1540,
		52364	=>	1541,
		52365	=>	1542,
		52366	=>	1543,
		52367	=>	1544,
		52368	=>	1545,
		52369	=>	1546,
		52370	=>	1547,
		52371	=>	1548,
		52372	=>	1549,
		52373	=>	1550,
		52374	=>	1551,
		52375	=>	1552,
		52376	=>	1553,
		52377	=>	1554,
		52378	=>	1555,
		52379	=>	1556,
		52380	=>	1557,
		52381	=>	1558,
		52382	=>	1559,
		52383	=>	1560,
		52384	=>	1561,
		52385	=>	1562,
		52386	=>	1562,
		52387	=>	1563,
		52388	=>	1564,
		52389	=>	1565,
		52390	=>	1566,
		52391	=>	1567,
		52392	=>	1568,
		52393	=>	1569,
		52394	=>	1570,
		52395	=>	1571,
		52396	=>	1572,
		52397	=>	1573,
		52398	=>	1574,
		52399	=>	1575,
		52400	=>	1576,
		52401	=>	1577,
		52402	=>	1578,
		52403	=>	1579,
		52404	=>	1580,
		52405	=>	1581,
		52406	=>	1582,
		52407	=>	1583,
		52408	=>	1584,
		52409	=>	1585,
		52410	=>	1586,
		52411	=>	1587,
		52412	=>	1587,
		52413	=>	1588,
		52414	=>	1589,
		52415	=>	1590,
		52416	=>	1591,
		52417	=>	1592,
		52418	=>	1593,
		52419	=>	1594,
		52420	=>	1595,
		52421	=>	1596,
		52422	=>	1597,
		52423	=>	1598,
		52424	=>	1599,
		52425	=>	1600,
		52426	=>	1601,
		52427	=>	1602,
		52428	=>	1603,
		52429	=>	1604,
		52430	=>	1605,
		52431	=>	1606,
		52432	=>	1607,
		52433	=>	1608,
		52434	=>	1609,
		52435	=>	1610,
		52436	=>	1611,
		52437	=>	1612,
		52438	=>	1613,
		52439	=>	1614,
		52440	=>	1615,
		52441	=>	1616,
		52442	=>	1617,
		52443	=>	1618,
		52444	=>	1619,
		52445	=>	1620,
		52446	=>	1620,
		52447	=>	1621,
		52448	=>	1622,
		52449	=>	1623,
		52450	=>	1624,
		52451	=>	1625,
		52452	=>	1626,
		52453	=>	1627,
		52454	=>	1628,
		52455	=>	1629,
		52456	=>	1630,
		52457	=>	1631,
		52458	=>	1632,
		52459	=>	1633,
		52460	=>	1634,
		52461	=>	1635,
		52462	=>	1636,
		52463	=>	1637,
		52464	=>	1638,
		52465	=>	1639,
		52466	=>	1640,
		52467	=>	1641,
		52468	=>	1642,
		52469	=>	1643,
		52470	=>	1644,
		52471	=>	1645,
		52472	=>	1646,
		52473	=>	1647,
		52474	=>	1648,
		52475	=>	1649,
		52476	=>	1650,
		52477	=>	1651,
		52478	=>	1652,
		52479	=>	1653,
		52480	=>	1654,
		52481	=>	1655,
		52482	=>	1656,
		52483	=>	1657,
		52484	=>	1658,
		52485	=>	1659,
		52486	=>	1660,
		52487	=>	1661,
		52488	=>	1662,
		52489	=>	1663,
		52490	=>	1664,
		52491	=>	1665,
		52492	=>	1666,
		52493	=>	1667,
		52494	=>	1668,
		52495	=>	1669,
		52496	=>	1670,
		52497	=>	1671,
		52498	=>	1672,
		52499	=>	1673,
		52500	=>	1674,
		52501	=>	1675,
		52502	=>	1676,
		52503	=>	1677,
		52504	=>	1678,
		52505	=>	1679,
		52506	=>	1680,
		52507	=>	1681,
		52508	=>	1682,
		52509	=>	1683,
		52510	=>	1684,
		52511	=>	1685,
		52512	=>	1686,
		52513	=>	1687,
		52514	=>	1688,
		52515	=>	1689,
		52516	=>	1689,
		52517	=>	1690,
		52518	=>	1691,
		52519	=>	1692,
		52520	=>	1693,
		52521	=>	1694,
		52522	=>	1695,
		52523	=>	1696,
		52524	=>	1697,
		52525	=>	1698,
		52526	=>	1699,
		52527	=>	1700,
		52528	=>	1701,
		52529	=>	1702,
		52530	=>	1703,
		52531	=>	1704,
		52532	=>	1705,
		52533	=>	1706,
		52534	=>	1707,
		52535	=>	1708,
		52536	=>	1709,
		52537	=>	1710,
		52538	=>	1711,
		52539	=>	1712,
		52540	=>	1713,
		52541	=>	1714,
		52542	=>	1715,
		52543	=>	1716,
		52544	=>	1717,
		52545	=>	1718,
		52546	=>	1719,
		52547	=>	1721,
		52548	=>	1722,
		52549	=>	1723,
		52550	=>	1724,
		52551	=>	1725,
		52552	=>	1726,
		52553	=>	1727,
		52554	=>	1728,
		52555	=>	1729,
		52556	=>	1730,
		52557	=>	1731,
		52558	=>	1732,
		52559	=>	1733,
		52560	=>	1734,
		52561	=>	1735,
		52562	=>	1736,
		52563	=>	1737,
		52564	=>	1738,
		52565	=>	1739,
		52566	=>	1740,
		52567	=>	1741,
		52568	=>	1742,
		52569	=>	1743,
		52570	=>	1744,
		52571	=>	1745,
		52572	=>	1746,
		52573	=>	1747,
		52574	=>	1748,
		52575	=>	1749,
		52576	=>	1750,
		52577	=>	1751,
		52578	=>	1752,
		52579	=>	1753,
		52580	=>	1754,
		52581	=>	1755,
		52582	=>	1756,
		52583	=>	1757,
		52584	=>	1758,
		52585	=>	1759,
		52586	=>	1760,
		52587	=>	1761,
		52588	=>	1762,
		52589	=>	1763,
		52590	=>	1764,
		52591	=>	1765,
		52592	=>	1766,
		52593	=>	1767,
		52594	=>	1768,
		52595	=>	1769,
		52596	=>	1770,
		52597	=>	1771,
		52598	=>	1772,
		52599	=>	1773,
		52600	=>	1774,
		52601	=>	1775,
		52602	=>	1776,
		52603	=>	1777,
		52604	=>	1778,
		52605	=>	1779,
		52606	=>	1780,
		52607	=>	1781,
		52608	=>	1782,
		52609	=>	1783,
		52610	=>	1784,
		52611	=>	1785,
		52612	=>	1786,
		52613	=>	1787,
		52614	=>	1788,
		52615	=>	1789,
		52616	=>	1790,
		52617	=>	1792,
		52618	=>	1793,
		52619	=>	1794,
		52620	=>	1795,
		52621	=>	1796,
		52622	=>	1797,
		52623	=>	1798,
		52624	=>	1799,
		52625	=>	1800,
		52626	=>	1801,
		52627	=>	1802,
		52628	=>	1803,
		52629	=>	1804,
		52630	=>	1805,
		52631	=>	1806,
		52632	=>	1807,
		52633	=>	1808,
		52634	=>	1809,
		52635	=>	1810,
		52636	=>	1811,
		52637	=>	1812,
		52638	=>	1813,
		52639	=>	1814,
		52640	=>	1815,
		52641	=>	1816,
		52642	=>	1817,
		52643	=>	1818,
		52644	=>	1819,
		52645	=>	1820,
		52646	=>	1821,
		52647	=>	1822,
		52648	=>	1823,
		52649	=>	1824,
		52650	=>	1825,
		52651	=>	1827,
		52652	=>	1828,
		52653	=>	1829,
		52654	=>	1830,
		52655	=>	1831,
		52656	=>	1832,
		52657	=>	1833,
		52658	=>	1834,
		52659	=>	1835,
		52660	=>	1836,
		52661	=>	1837,
		52662	=>	1838,
		52663	=>	1839,
		52664	=>	1840,
		52665	=>	1841,
		52666	=>	1842,
		52667	=>	1843,
		52668	=>	1844,
		52669	=>	1845,
		52670	=>	1846,
		52671	=>	1847,
		52672	=>	1848,
		52673	=>	1849,
		52674	=>	1850,
		52675	=>	1851,
		52676	=>	1852,
		52677	=>	1854,
		52678	=>	1855,
		52679	=>	1856,
		52680	=>	1857,
		52681	=>	1858,
		52682	=>	1859,
		52683	=>	1860,
		52684	=>	1861,
		52685	=>	1862,
		52686	=>	1863,
		52687	=>	1864,
		52688	=>	1865,
		52689	=>	1866,
		52690	=>	1867,
		52691	=>	1868,
		52692	=>	1869,
		52693	=>	1870,
		52694	=>	1871,
		52695	=>	1872,
		52696	=>	1873,
		52697	=>	1874,
		52698	=>	1875,
		52699	=>	1876,
		52700	=>	1878,
		52701	=>	1879,
		52702	=>	1880,
		52703	=>	1881,
		52704	=>	1882,
		52705	=>	1883,
		52706	=>	1884,
		52707	=>	1885,
		52708	=>	1886,
		52709	=>	1887,
		52710	=>	1888,
		52711	=>	1889,
		52712	=>	1890,
		52713	=>	1891,
		52714	=>	1892,
		52715	=>	1893,
		52716	=>	1894,
		52717	=>	1895,
		52718	=>	1896,
		52719	=>	1898,
		52720	=>	1899,
		52721	=>	1900,
		52722	=>	1901,
		52723	=>	1902,
		52724	=>	1903,
		52725	=>	1904,
		52726	=>	1905,
		52727	=>	1906,
		52728	=>	1907,
		52729	=>	1908,
		52730	=>	1909,
		52731	=>	1910,
		52732	=>	1911,
		52733	=>	1912,
		52734	=>	1913,
		52735	=>	1914,
		52736	=>	1915,
		52737	=>	1917,
		52738	=>	1918,
		52739	=>	1919,
		52740	=>	1920,
		52741	=>	1921,
		52742	=>	1922,
		52743	=>	1923,
		52744	=>	1924,
		52745	=>	1925,
		52746	=>	1926,
		52747	=>	1927,
		52748	=>	1928,
		52749	=>	1929,
		52750	=>	1930,
		52751	=>	1931,
		52752	=>	1932,
		52753	=>	1933,
		52754	=>	1935,
		52755	=>	1936,
		52756	=>	1937,
		52757	=>	1938,
		52758	=>	1939,
		52759	=>	1940,
		52760	=>	1941,
		52761	=>	1942,
		52762	=>	1943,
		52763	=>	1944,
		52764	=>	1945,
		52765	=>	1946,
		52766	=>	1947,
		52767	=>	1948,
		52768	=>	1949,
		52769	=>	1951,
		52770	=>	1952,
		52771	=>	1953,
		52772	=>	1954,
		52773	=>	1955,
		52774	=>	1956,
		52775	=>	1957,
		52776	=>	1958,
		52777	=>	1959,
		52778	=>	1960,
		52779	=>	1961,
		52780	=>	1962,
		52781	=>	1963,
		52782	=>	1964,
		52783	=>	1966,
		52784	=>	1967,
		52785	=>	1968,
		52786	=>	1969,
		52787	=>	1970,
		52788	=>	1971,
		52789	=>	1972,
		52790	=>	1973,
		52791	=>	1974,
		52792	=>	1975,
		52793	=>	1976,
		52794	=>	1977,
		52795	=>	1978,
		52796	=>	1979,
		52797	=>	1981,
		52798	=>	1982,
		52799	=>	1983,
		52800	=>	1984,
		52801	=>	1985,
		52802	=>	1986,
		52803	=>	1987,
		52804	=>	1988,
		52805	=>	1989,
		52806	=>	1990,
		52807	=>	1991,
		52808	=>	1992,
		52809	=>	1993,
		52810	=>	1995,
		52811	=>	1996,
		52812	=>	1997,
		52813	=>	1998,
		52814	=>	1999,
		52815	=>	2000,
		52816	=>	2001,
		52817	=>	2002,
		52818	=>	2003,
		52819	=>	2004,
		52820	=>	2005,
		52821	=>	2006,
		52822	=>	2008,
		52823	=>	2009,
		52824	=>	2010,
		52825	=>	2011,
		52826	=>	2012,
		52827	=>	2013,
		52828	=>	2014,
		52829	=>	2015,
		52830	=>	2016,
		52831	=>	2017,
		52832	=>	2018,
		52833	=>	2019,
		52834	=>	2021,
		52835	=>	2022,
		52836	=>	2023,
		52837	=>	2024,
		52838	=>	2025,
		52839	=>	2026,
		52840	=>	2027,
		52841	=>	2028,
		52842	=>	2029,
		52843	=>	2030,
		52844	=>	2031,
		52845	=>	2032,
		52846	=>	2034,
		52847	=>	2035,
		52848	=>	2036,
		52849	=>	2037,
		52850	=>	2038,
		52851	=>	2039,
		52852	=>	2040,
		52853	=>	2041,
		52854	=>	2042,
		52855	=>	2043,
		52856	=>	2044,
		52857	=>	2046,
		52858	=>	2047,
		52859	=>	2048,
		52860	=>	2049,
		52861	=>	2050,
		52862	=>	2051,
		52863	=>	2052,
		52864	=>	2053,
		52865	=>	2054,
		52866	=>	2055,
		52867	=>	2057,
		52868	=>	2058,
		52869	=>	2059,
		52870	=>	2060,
		52871	=>	2061,
		52872	=>	2062,
		52873	=>	2063,
		52874	=>	2064,
		52875	=>	2065,
		52876	=>	2066,
		52877	=>	2067,
		52878	=>	2069,
		52879	=>	2070,
		52880	=>	2071,
		52881	=>	2072,
		52882	=>	2073,
		52883	=>	2074,
		52884	=>	2075,
		52885	=>	2076,
		52886	=>	2077,
		52887	=>	2078,
		52888	=>	2080,
		52889	=>	2081,
		52890	=>	2082,
		52891	=>	2083,
		52892	=>	2084,
		52893	=>	2085,
		52894	=>	2086,
		52895	=>	2087,
		52896	=>	2088,
		52897	=>	2090,
		52898	=>	2091,
		52899	=>	2092,
		52900	=>	2093,
		52901	=>	2094,
		52902	=>	2095,
		52903	=>	2096,
		52904	=>	2097,
		52905	=>	2098,
		52906	=>	2099,
		52907	=>	2101,
		52908	=>	2102,
		52909	=>	2103,
		52910	=>	2104,
		52911	=>	2105,
		52912	=>	2106,
		52913	=>	2107,
		52914	=>	2108,
		52915	=>	2109,
		52916	=>	2111,
		52917	=>	2112,
		52918	=>	2113,
		52919	=>	2114,
		52920	=>	2115,
		52921	=>	2116,
		52922	=>	2117,
		52923	=>	2118,
		52924	=>	2119,
		52925	=>	2121,
		52926	=>	2122,
		52927	=>	2123,
		52928	=>	2124,
		52929	=>	2125,
		52930	=>	2126,
		52931	=>	2127,
		52932	=>	2128,
		52933	=>	2129,
		52934	=>	2131,
		52935	=>	2132,
		52936	=>	2133,
		52937	=>	2134,
		52938	=>	2135,
		52939	=>	2136,
		52940	=>	2137,
		52941	=>	2138,
		52942	=>	2139,
		52943	=>	2141,
		52944	=>	2142,
		52945	=>	2143,
		52946	=>	2144,
		52947	=>	2145,
		52948	=>	2146,
		52949	=>	2147,
		52950	=>	2148,
		52951	=>	2150,
		52952	=>	2151,
		52953	=>	2152,
		52954	=>	2153,
		52955	=>	2154,
		52956	=>	2155,
		52957	=>	2156,
		52958	=>	2157,
		52959	=>	2159,
		52960	=>	2160,
		52961	=>	2161,
		52962	=>	2162,
		52963	=>	2163,
		52964	=>	2164,
		52965	=>	2165,
		52966	=>	2166,
		52967	=>	2167,
		52968	=>	2169,
		52969	=>	2170,
		52970	=>	2171,
		52971	=>	2172,
		52972	=>	2173,
		52973	=>	2174,
		52974	=>	2175,
		52975	=>	2176,
		52976	=>	2178,
		52977	=>	2179,
		52978	=>	2180,
		52979	=>	2181,
		52980	=>	2182,
		52981	=>	2183,
		52982	=>	2184,
		52983	=>	2185,
		52984	=>	2187,
		52985	=>	2188,
		52986	=>	2189,
		52987	=>	2190,
		52988	=>	2191,
		52989	=>	2192,
		52990	=>	2193,
		52991	=>	2195,
		52992	=>	2196,
		52993	=>	2197,
		52994	=>	2198,
		52995	=>	2199,
		52996	=>	2200,
		52997	=>	2201,
		52998	=>	2202,
		52999	=>	2204,
		53000	=>	2205,
		53001	=>	2206,
		53002	=>	2207,
		53003	=>	2208,
		53004	=>	2209,
		53005	=>	2210,
		53006	=>	2212,
		53007	=>	2213,
		53008	=>	2214,
		53009	=>	2215,
		53010	=>	2216,
		53011	=>	2217,
		53012	=>	2218,
		53013	=>	2219,
		53014	=>	2221,
		53015	=>	2222,
		53016	=>	2223,
		53017	=>	2224,
		53018	=>	2225,
		53019	=>	2226,
		53020	=>	2227,
		53021	=>	2229,
		53022	=>	2230,
		53023	=>	2231,
		53024	=>	2232,
		53025	=>	2233,
		53026	=>	2234,
		53027	=>	2235,
		53028	=>	2237,
		53029	=>	2238,
		53030	=>	2239,
		53031	=>	2240,
		53032	=>	2241,
		53033	=>	2242,
		53034	=>	2243,
		53035	=>	2245,
		53036	=>	2246,
		53037	=>	2247,
		53038	=>	2248,
		53039	=>	2249,
		53040	=>	2250,
		53041	=>	2251,
		53042	=>	2253,
		53043	=>	2254,
		53044	=>	2255,
		53045	=>	2256,
		53046	=>	2257,
		53047	=>	2258,
		53048	=>	2259,
		53049	=>	2261,
		53050	=>	2262,
		53051	=>	2263,
		53052	=>	2264,
		53053	=>	2265,
		53054	=>	2266,
		53055	=>	2267,
		53056	=>	2269,
		53057	=>	2270,
		53058	=>	2271,
		53059	=>	2272,
		53060	=>	2273,
		53061	=>	2274,
		53062	=>	2275,
		53063	=>	2277,
		53064	=>	2278,
		53065	=>	2279,
		53066	=>	2280,
		53067	=>	2281,
		53068	=>	2282,
		53069	=>	2284,
		53070	=>	2285,
		53071	=>	2286,
		53072	=>	2287,
		53073	=>	2288,
		53074	=>	2289,
		53075	=>	2290,
		53076	=>	2292,
		53077	=>	2293,
		53078	=>	2294,
		53079	=>	2295,
		53080	=>	2296,
		53081	=>	2297,
		53082	=>	2299,
		53083	=>	2300,
		53084	=>	2301,
		53085	=>	2302,
		53086	=>	2303,
		53087	=>	2304,
		53088	=>	2305,
		53089	=>	2307,
		53090	=>	2308,
		53091	=>	2309,
		53092	=>	2310,
		53093	=>	2311,
		53094	=>	2312,
		53095	=>	2314,
		53096	=>	2315,
		53097	=>	2316,
		53098	=>	2317,
		53099	=>	2318,
		53100	=>	2319,
		53101	=>	2321,
		53102	=>	2322,
		53103	=>	2323,
		53104	=>	2324,
		53105	=>	2325,
		53106	=>	2326,
		53107	=>	2328,
		53108	=>	2329,
		53109	=>	2330,
		53110	=>	2331,
		53111	=>	2332,
		53112	=>	2333,
		53113	=>	2335,
		53114	=>	2336,
		53115	=>	2337,
		53116	=>	2338,
		53117	=>	2339,
		53118	=>	2340,
		53119	=>	2342,
		53120	=>	2343,
		53121	=>	2344,
		53122	=>	2345,
		53123	=>	2346,
		53124	=>	2347,
		53125	=>	2349,
		53126	=>	2350,
		53127	=>	2351,
		53128	=>	2352,
		53129	=>	2353,
		53130	=>	2354,
		53131	=>	2356,
		53132	=>	2357,
		53133	=>	2358,
		53134	=>	2359,
		53135	=>	2360,
		53136	=>	2361,
		53137	=>	2363,
		53138	=>	2364,
		53139	=>	2365,
		53140	=>	2366,
		53141	=>	2367,
		53142	=>	2368,
		53143	=>	2370,
		53144	=>	2371,
		53145	=>	2372,
		53146	=>	2373,
		53147	=>	2374,
		53148	=>	2375,
		53149	=>	2377,
		53150	=>	2378,
		53151	=>	2379,
		53152	=>	2380,
		53153	=>	2381,
		53154	=>	2382,
		53155	=>	2384,
		53156	=>	2385,
		53157	=>	2386,
		53158	=>	2387,
		53159	=>	2388,
		53160	=>	2390,
		53161	=>	2391,
		53162	=>	2392,
		53163	=>	2393,
		53164	=>	2394,
		53165	=>	2395,
		53166	=>	2397,
		53167	=>	2398,
		53168	=>	2399,
		53169	=>	2400,
		53170	=>	2401,
		53171	=>	2403,
		53172	=>	2404,
		53173	=>	2405,
		53174	=>	2406,
		53175	=>	2407,
		53176	=>	2408,
		53177	=>	2410,
		53178	=>	2411,
		53179	=>	2412,
		53180	=>	2413,
		53181	=>	2414,
		53182	=>	2416,
		53183	=>	2417,
		53184	=>	2418,
		53185	=>	2419,
		53186	=>	2420,
		53187	=>	2421,
		53188	=>	2423,
		53189	=>	2424,
		53190	=>	2425,
		53191	=>	2426,
		53192	=>	2427,
		53193	=>	2429,
		53194	=>	2430,
		53195	=>	2431,
		53196	=>	2432,
		53197	=>	2433,
		53198	=>	2435,
		53199	=>	2436,
		53200	=>	2437,
		53201	=>	2438,
		53202	=>	2439,
		53203	=>	2440,
		53204	=>	2442,
		53205	=>	2443,
		53206	=>	2444,
		53207	=>	2445,
		53208	=>	2446,
		53209	=>	2448,
		53210	=>	2449,
		53211	=>	2450,
		53212	=>	2451,
		53213	=>	2452,
		53214	=>	2454,
		53215	=>	2455,
		53216	=>	2456,
		53217	=>	2457,
		53218	=>	2458,
		53219	=>	2460,
		53220	=>	2461,
		53221	=>	2462,
		53222	=>	2463,
		53223	=>	2464,
		53224	=>	2466,
		53225	=>	2467,
		53226	=>	2468,
		53227	=>	2469,
		53228	=>	2470,
		53229	=>	2471,
		53230	=>	2473,
		53231	=>	2474,
		53232	=>	2475,
		53233	=>	2476,
		53234	=>	2477,
		53235	=>	2479,
		53236	=>	2480,
		53237	=>	2481,
		53238	=>	2482,
		53239	=>	2483,
		53240	=>	2485,
		53241	=>	2486,
		53242	=>	2487,
		53243	=>	2488,
		53244	=>	2489,
		53245	=>	2491,
		53246	=>	2492,
		53247	=>	2493,
		53248	=>	2494,
		53249	=>	2495,
		53250	=>	2497,
		53251	=>	2498,
		53252	=>	2499,
		53253	=>	2500,
		53254	=>	2501,
		53255	=>	2503,
		53256	=>	2504,
		53257	=>	2505,
		53258	=>	2506,
		53259	=>	2508,
		53260	=>	2509,
		53261	=>	2510,
		53262	=>	2511,
		53263	=>	2512,
		53264	=>	2514,
		53265	=>	2515,
		53266	=>	2516,
		53267	=>	2517,
		53268	=>	2518,
		53269	=>	2520,
		53270	=>	2521,
		53271	=>	2522,
		53272	=>	2523,
		53273	=>	2524,
		53274	=>	2526,
		53275	=>	2527,
		53276	=>	2528,
		53277	=>	2529,
		53278	=>	2530,
		53279	=>	2532,
		53280	=>	2533,
		53281	=>	2534,
		53282	=>	2535,
		53283	=>	2537,
		53284	=>	2538,
		53285	=>	2539,
		53286	=>	2540,
		53287	=>	2541,
		53288	=>	2543,
		53289	=>	2544,
		53290	=>	2545,
		53291	=>	2546,
		53292	=>	2547,
		53293	=>	2549,
		53294	=>	2550,
		53295	=>	2551,
		53296	=>	2552,
		53297	=>	2554,
		53298	=>	2555,
		53299	=>	2556,
		53300	=>	2557,
		53301	=>	2558,
		53302	=>	2560,
		53303	=>	2561,
		53304	=>	2562,
		53305	=>	2563,
		53306	=>	2564,
		53307	=>	2566,
		53308	=>	2567,
		53309	=>	2568,
		53310	=>	2569,
		53311	=>	2571,
		53312	=>	2572,
		53313	=>	2573,
		53314	=>	2574,
		53315	=>	2575,
		53316	=>	2577,
		53317	=>	2578,
		53318	=>	2579,
		53319	=>	2580,
		53320	=>	2582,
		53321	=>	2583,
		53322	=>	2584,
		53323	=>	2585,
		53324	=>	2586,
		53325	=>	2588,
		53326	=>	2589,
		53327	=>	2590,
		53328	=>	2591,
		53329	=>	2593,
		53330	=>	2594,
		53331	=>	2595,
		53332	=>	2596,
		53333	=>	2597,
		53334	=>	2599,
		53335	=>	2600,
		53336	=>	2601,
		53337	=>	2602,
		53338	=>	2604,
		53339	=>	2605,
		53340	=>	2606,
		53341	=>	2607,
		53342	=>	2609,
		53343	=>	2610,
		53344	=>	2611,
		53345	=>	2612,
		53346	=>	2613,
		53347	=>	2615,
		53348	=>	2616,
		53349	=>	2617,
		53350	=>	2618,
		53351	=>	2620,
		53352	=>	2621,
		53353	=>	2622,
		53354	=>	2623,
		53355	=>	2625,
		53356	=>	2626,
		53357	=>	2627,
		53358	=>	2628,
		53359	=>	2629,
		53360	=>	2631,
		53361	=>	2632,
		53362	=>	2633,
		53363	=>	2634,
		53364	=>	2636,
		53365	=>	2637,
		53366	=>	2638,
		53367	=>	2639,
		53368	=>	2641,
		53369	=>	2642,
		53370	=>	2643,
		53371	=>	2644,
		53372	=>	2645,
		53373	=>	2647,
		53374	=>	2648,
		53375	=>	2649,
		53376	=>	2650,
		53377	=>	2652,
		53378	=>	2653,
		53379	=>	2654,
		53380	=>	2655,
		53381	=>	2657,
		53382	=>	2658,
		53383	=>	2659,
		53384	=>	2660,
		53385	=>	2662,
		53386	=>	2663,
		53387	=>	2664,
		53388	=>	2665,
		53389	=>	2667,
		53390	=>	2668,
		53391	=>	2669,
		53392	=>	2670,
		53393	=>	2672,
		53394	=>	2673,
		53395	=>	2674,
		53396	=>	2675,
		53397	=>	2676,
		53398	=>	2678,
		53399	=>	2679,
		53400	=>	2680,
		53401	=>	2681,
		53402	=>	2683,
		53403	=>	2684,
		53404	=>	2685,
		53405	=>	2686,
		53406	=>	2688,
		53407	=>	2689,
		53408	=>	2690,
		53409	=>	2691,
		53410	=>	2693,
		53411	=>	2694,
		53412	=>	2695,
		53413	=>	2696,
		53414	=>	2698,
		53415	=>	2699,
		53416	=>	2700,
		53417	=>	2701,
		53418	=>	2703,
		53419	=>	2704,
		53420	=>	2705,
		53421	=>	2706,
		53422	=>	2708,
		53423	=>	2709,
		53424	=>	2710,
		53425	=>	2711,
		53426	=>	2713,
		53427	=>	2714,
		53428	=>	2715,
		53429	=>	2716,
		53430	=>	2718,
		53431	=>	2719,
		53432	=>	2720,
		53433	=>	2721,
		53434	=>	2723,
		53435	=>	2724,
		53436	=>	2725,
		53437	=>	2726,
		53438	=>	2728,
		53439	=>	2729,
		53440	=>	2730,
		53441	=>	2731,
		53442	=>	2733,
		53443	=>	2734,
		53444	=>	2735,
		53445	=>	2736,
		53446	=>	2738,
		53447	=>	2739,
		53448	=>	2740,
		53449	=>	2742,
		53450	=>	2743,
		53451	=>	2744,
		53452	=>	2745,
		53453	=>	2747,
		53454	=>	2748,
		53455	=>	2749,
		53456	=>	2750,
		53457	=>	2752,
		53458	=>	2753,
		53459	=>	2754,
		53460	=>	2755,
		53461	=>	2757,
		53462	=>	2758,
		53463	=>	2759,
		53464	=>	2760,
		53465	=>	2762,
		53466	=>	2763,
		53467	=>	2764,
		53468	=>	2765,
		53469	=>	2767,
		53470	=>	2768,
		53471	=>	2769,
		53472	=>	2771,
		53473	=>	2772,
		53474	=>	2773,
		53475	=>	2774,
		53476	=>	2776,
		53477	=>	2777,
		53478	=>	2778,
		53479	=>	2779,
		53480	=>	2781,
		53481	=>	2782,
		53482	=>	2783,
		53483	=>	2784,
		53484	=>	2786,
		53485	=>	2787,
		53486	=>	2788,
		53487	=>	2790,
		53488	=>	2791,
		53489	=>	2792,
		53490	=>	2793,
		53491	=>	2795,
		53492	=>	2796,
		53493	=>	2797,
		53494	=>	2798,
		53495	=>	2800,
		53496	=>	2801,
		53497	=>	2802,
		53498	=>	2803,
		53499	=>	2805,
		53500	=>	2806,
		53501	=>	2807,
		53502	=>	2809,
		53503	=>	2810,
		53504	=>	2811,
		53505	=>	2812,
		53506	=>	2814,
		53507	=>	2815,
		53508	=>	2816,
		53509	=>	2818,
		53510	=>	2819,
		53511	=>	2820,
		53512	=>	2821,
		53513	=>	2823,
		53514	=>	2824,
		53515	=>	2825,
		53516	=>	2826,
		53517	=>	2828,
		53518	=>	2829,
		53519	=>	2830,
		53520	=>	2832,
		53521	=>	2833,
		53522	=>	2834,
		53523	=>	2835,
		53524	=>	2837,
		53525	=>	2838,
		53526	=>	2839,
		53527	=>	2840,
		53528	=>	2842,
		53529	=>	2843,
		53530	=>	2844,
		53531	=>	2846,
		53532	=>	2847,
		53533	=>	2848,
		53534	=>	2849,
		53535	=>	2851,
		53536	=>	2852,
		53537	=>	2853,
		53538	=>	2855,
		53539	=>	2856,
		53540	=>	2857,
		53541	=>	2858,
		53542	=>	2860,
		53543	=>	2861,
		53544	=>	2862,
		53545	=>	2864,
		53546	=>	2865,
		53547	=>	2866,
		53548	=>	2867,
		53549	=>	2869,
		53550	=>	2870,
		53551	=>	2871,
		53552	=>	2873,
		53553	=>	2874,
		53554	=>	2875,
		53555	=>	2876,
		53556	=>	2878,
		53557	=>	2879,
		53558	=>	2880,
		53559	=>	2882,
		53560	=>	2883,
		53561	=>	2884,
		53562	=>	2885,
		53563	=>	2887,
		53564	=>	2888,
		53565	=>	2889,
		53566	=>	2891,
		53567	=>	2892,
		53568	=>	2893,
		53569	=>	2894,
		53570	=>	2896,
		53571	=>	2897,
		53572	=>	2898,
		53573	=>	2900,
		53574	=>	2901,
		53575	=>	2902,
		53576	=>	2904,
		53577	=>	2905,
		53578	=>	2906,
		53579	=>	2907,
		53580	=>	2909,
		53581	=>	2910,
		53582	=>	2911,
		53583	=>	2913,
		53584	=>	2914,
		53585	=>	2915,
		53586	=>	2916,
		53587	=>	2918,
		53588	=>	2919,
		53589	=>	2920,
		53590	=>	2922,
		53591	=>	2923,
		53592	=>	2924,
		53593	=>	2926,
		53594	=>	2927,
		53595	=>	2928,
		53596	=>	2929,
		53597	=>	2931,
		53598	=>	2932,
		53599	=>	2933,
		53600	=>	2935,
		53601	=>	2936,
		53602	=>	2937,
		53603	=>	2939,
		53604	=>	2940,
		53605	=>	2941,
		53606	=>	2942,
		53607	=>	2944,
		53608	=>	2945,
		53609	=>	2946,
		53610	=>	2948,
		53611	=>	2949,
		53612	=>	2950,
		53613	=>	2952,
		53614	=>	2953,
		53615	=>	2954,
		53616	=>	2955,
		53617	=>	2957,
		53618	=>	2958,
		53619	=>	2959,
		53620	=>	2961,
		53621	=>	2962,
		53622	=>	2963,
		53623	=>	2965,
		53624	=>	2966,
		53625	=>	2967,
		53626	=>	2968,
		53627	=>	2970,
		53628	=>	2971,
		53629	=>	2972,
		53630	=>	2974,
		53631	=>	2975,
		53632	=>	2976,
		53633	=>	2978,
		53634	=>	2979,
		53635	=>	2980,
		53636	=>	2982,
		53637	=>	2983,
		53638	=>	2984,
		53639	=>	2986,
		53640	=>	2987,
		53641	=>	2988,
		53642	=>	2989,
		53643	=>	2991,
		53644	=>	2992,
		53645	=>	2993,
		53646	=>	2995,
		53647	=>	2996,
		53648	=>	2997,
		53649	=>	2999,
		53650	=>	3000,
		53651	=>	3001,
		53652	=>	3003,
		53653	=>	3004,
		53654	=>	3005,
		53655	=>	3006,
		53656	=>	3008,
		53657	=>	3009,
		53658	=>	3010,
		53659	=>	3012,
		53660	=>	3013,
		53661	=>	3014,
		53662	=>	3016,
		53663	=>	3017,
		53664	=>	3018,
		53665	=>	3020,
		53666	=>	3021,
		53667	=>	3022,
		53668	=>	3024,
		53669	=>	3025,
		53670	=>	3026,
		53671	=>	3028,
		53672	=>	3029,
		53673	=>	3030,
		53674	=>	3032,
		53675	=>	3033,
		53676	=>	3034,
		53677	=>	3035,
		53678	=>	3037,
		53679	=>	3038,
		53680	=>	3039,
		53681	=>	3041,
		53682	=>	3042,
		53683	=>	3043,
		53684	=>	3045,
		53685	=>	3046,
		53686	=>	3047,
		53687	=>	3049,
		53688	=>	3050,
		53689	=>	3051,
		53690	=>	3053,
		53691	=>	3054,
		53692	=>	3055,
		53693	=>	3057,
		53694	=>	3058,
		53695	=>	3059,
		53696	=>	3061,
		53697	=>	3062,
		53698	=>	3063,
		53699	=>	3065,
		53700	=>	3066,
		53701	=>	3067,
		53702	=>	3069,
		53703	=>	3070,
		53704	=>	3071,
		53705	=>	3073,
		53706	=>	3074,
		53707	=>	3075,
		53708	=>	3077,
		53709	=>	3078,
		53710	=>	3079,
		53711	=>	3081,
		53712	=>	3082,
		53713	=>	3083,
		53714	=>	3085,
		53715	=>	3086,
		53716	=>	3087,
		53717	=>	3089,
		53718	=>	3090,
		53719	=>	3091,
		53720	=>	3093,
		53721	=>	3094,
		53722	=>	3095,
		53723	=>	3097,
		53724	=>	3098,
		53725	=>	3099,
		53726	=>	3101,
		53727	=>	3102,
		53728	=>	3103,
		53729	=>	3105,
		53730	=>	3106,
		53731	=>	3107,
		53732	=>	3109,
		53733	=>	3110,
		53734	=>	3111,
		53735	=>	3113,
		53736	=>	3114,
		53737	=>	3115,
		53738	=>	3117,
		53739	=>	3118,
		53740	=>	3119,
		53741	=>	3121,
		53742	=>	3122,
		53743	=>	3123,
		53744	=>	3125,
		53745	=>	3126,
		53746	=>	3127,
		53747	=>	3129,
		53748	=>	3130,
		53749	=>	3131,
		53750	=>	3133,
		53751	=>	3134,
		53752	=>	3135,
		53753	=>	3137,
		53754	=>	3138,
		53755	=>	3139,
		53756	=>	3141,
		53757	=>	3142,
		53758	=>	3143,
		53759	=>	3145,
		53760	=>	3146,
		53761	=>	3147,
		53762	=>	3149,
		53763	=>	3150,
		53764	=>	3151,
		53765	=>	3153,
		53766	=>	3154,
		53767	=>	3155,
		53768	=>	3157,
		53769	=>	3158,
		53770	=>	3159,
		53771	=>	3161,
		53772	=>	3162,
		53773	=>	3164,
		53774	=>	3165,
		53775	=>	3166,
		53776	=>	3168,
		53777	=>	3169,
		53778	=>	3170,
		53779	=>	3172,
		53780	=>	3173,
		53781	=>	3174,
		53782	=>	3176,
		53783	=>	3177,
		53784	=>	3178,
		53785	=>	3180,
		53786	=>	3181,
		53787	=>	3182,
		53788	=>	3184,
		53789	=>	3185,
		53790	=>	3186,
		53791	=>	3188,
		53792	=>	3189,
		53793	=>	3191,
		53794	=>	3192,
		53795	=>	3193,
		53796	=>	3195,
		53797	=>	3196,
		53798	=>	3197,
		53799	=>	3199,
		53800	=>	3200,
		53801	=>	3201,
		53802	=>	3203,
		53803	=>	3204,
		53804	=>	3205,
		53805	=>	3207,
		53806	=>	3208,
		53807	=>	3209,
		53808	=>	3211,
		53809	=>	3212,
		53810	=>	3214,
		53811	=>	3215,
		53812	=>	3216,
		53813	=>	3218,
		53814	=>	3219,
		53815	=>	3220,
		53816	=>	3222,
		53817	=>	3223,
		53818	=>	3224,
		53819	=>	3226,
		53820	=>	3227,
		53821	=>	3228,
		53822	=>	3230,
		53823	=>	3231,
		53824	=>	3233,
		53825	=>	3234,
		53826	=>	3235,
		53827	=>	3237,
		53828	=>	3238,
		53829	=>	3239,
		53830	=>	3241,
		53831	=>	3242,
		53832	=>	3243,
		53833	=>	3245,
		53834	=>	3246,
		53835	=>	3248,
		53836	=>	3249,
		53837	=>	3250,
		53838	=>	3252,
		53839	=>	3253,
		53840	=>	3254,
		53841	=>	3256,
		53842	=>	3257,
		53843	=>	3258,
		53844	=>	3260,
		53845	=>	3261,
		53846	=>	3263,
		53847	=>	3264,
		53848	=>	3265,
		53849	=>	3267,
		53850	=>	3268,
		53851	=>	3269,
		53852	=>	3271,
		53853	=>	3272,
		53854	=>	3273,
		53855	=>	3275,
		53856	=>	3276,
		53857	=>	3278,
		53858	=>	3279,
		53859	=>	3280,
		53860	=>	3282,
		53861	=>	3283,
		53862	=>	3284,
		53863	=>	3286,
		53864	=>	3287,
		53865	=>	3289,
		53866	=>	3290,
		53867	=>	3291,
		53868	=>	3293,
		53869	=>	3294,
		53870	=>	3295,
		53871	=>	3297,
		53872	=>	3298,
		53873	=>	3300,
		53874	=>	3301,
		53875	=>	3302,
		53876	=>	3304,
		53877	=>	3305,
		53878	=>	3306,
		53879	=>	3308,
		53880	=>	3309,
		53881	=>	3311,
		53882	=>	3312,
		53883	=>	3313,
		53884	=>	3315,
		53885	=>	3316,
		53886	=>	3317,
		53887	=>	3319,
		53888	=>	3320,
		53889	=>	3322,
		53890	=>	3323,
		53891	=>	3324,
		53892	=>	3326,
		53893	=>	3327,
		53894	=>	3328,
		53895	=>	3330,
		53896	=>	3331,
		53897	=>	3333,
		53898	=>	3334,
		53899	=>	3335,
		53900	=>	3337,
		53901	=>	3338,
		53902	=>	3340,
		53903	=>	3341,
		53904	=>	3342,
		53905	=>	3344,
		53906	=>	3345,
		53907	=>	3346,
		53908	=>	3348,
		53909	=>	3349,
		53910	=>	3351,
		53911	=>	3352,
		53912	=>	3353,
		53913	=>	3355,
		53914	=>	3356,
		53915	=>	3357,
		53916	=>	3359,
		53917	=>	3360,
		53918	=>	3362,
		53919	=>	3363,
		53920	=>	3364,
		53921	=>	3366,
		53922	=>	3367,
		53923	=>	3369,
		53924	=>	3370,
		53925	=>	3371,
		53926	=>	3373,
		53927	=>	3374,
		53928	=>	3376,
		53929	=>	3377,
		53930	=>	3378,
		53931	=>	3380,
		53932	=>	3381,
		53933	=>	3382,
		53934	=>	3384,
		53935	=>	3385,
		53936	=>	3387,
		53937	=>	3388,
		53938	=>	3389,
		53939	=>	3391,
		53940	=>	3392,
		53941	=>	3394,
		53942	=>	3395,
		53943	=>	3396,
		53944	=>	3398,
		53945	=>	3399,
		53946	=>	3401,
		53947	=>	3402,
		53948	=>	3403,
		53949	=>	3405,
		53950	=>	3406,
		53951	=>	3408,
		53952	=>	3409,
		53953	=>	3410,
		53954	=>	3412,
		53955	=>	3413,
		53956	=>	3415,
		53957	=>	3416,
		53958	=>	3417,
		53959	=>	3419,
		53960	=>	3420,
		53961	=>	3421,
		53962	=>	3423,
		53963	=>	3424,
		53964	=>	3426,
		53965	=>	3427,
		53966	=>	3428,
		53967	=>	3430,
		53968	=>	3431,
		53969	=>	3433,
		53970	=>	3434,
		53971	=>	3435,
		53972	=>	3437,
		53973	=>	3438,
		53974	=>	3440,
		53975	=>	3441,
		53976	=>	3442,
		53977	=>	3444,
		53978	=>	3445,
		53979	=>	3447,
		53980	=>	3448,
		53981	=>	3450,
		53982	=>	3451,
		53983	=>	3452,
		53984	=>	3454,
		53985	=>	3455,
		53986	=>	3457,
		53987	=>	3458,
		53988	=>	3459,
		53989	=>	3461,
		53990	=>	3462,
		53991	=>	3464,
		53992	=>	3465,
		53993	=>	3466,
		53994	=>	3468,
		53995	=>	3469,
		53996	=>	3471,
		53997	=>	3472,
		53998	=>	3473,
		53999	=>	3475,
		54000	=>	3476,
		54001	=>	3478,
		54002	=>	3479,
		54003	=>	3480,
		54004	=>	3482,
		54005	=>	3483,
		54006	=>	3485,
		54007	=>	3486,
		54008	=>	3487,
		54009	=>	3489,
		54010	=>	3490,
		54011	=>	3492,
		54012	=>	3493,
		54013	=>	3495,
		54014	=>	3496,
		54015	=>	3497,
		54016	=>	3499,
		54017	=>	3500,
		54018	=>	3502,
		54019	=>	3503,
		54020	=>	3504,
		54021	=>	3506,
		54022	=>	3507,
		54023	=>	3509,
		54024	=>	3510,
		54025	=>	3511,
		54026	=>	3513,
		54027	=>	3514,
		54028	=>	3516,
		54029	=>	3517,
		54030	=>	3519,
		54031	=>	3520,
		54032	=>	3521,
		54033	=>	3523,
		54034	=>	3524,
		54035	=>	3526,
		54036	=>	3527,
		54037	=>	3528,
		54038	=>	3530,
		54039	=>	3531,
		54040	=>	3533,
		54041	=>	3534,
		54042	=>	3536,
		54043	=>	3537,
		54044	=>	3538,
		54045	=>	3540,
		54046	=>	3541,
		54047	=>	3543,
		54048	=>	3544,
		54049	=>	3546,
		54050	=>	3547,
		54051	=>	3548,
		54052	=>	3550,
		54053	=>	3551,
		54054	=>	3553,
		54055	=>	3554,
		54056	=>	3555,
		54057	=>	3557,
		54058	=>	3558,
		54059	=>	3560,
		54060	=>	3561,
		54061	=>	3563,
		54062	=>	3564,
		54063	=>	3565,
		54064	=>	3567,
		54065	=>	3568,
		54066	=>	3570,
		54067	=>	3571,
		54068	=>	3573,
		54069	=>	3574,
		54070	=>	3575,
		54071	=>	3577,
		54072	=>	3578,
		54073	=>	3580,
		54074	=>	3581,
		54075	=>	3583,
		54076	=>	3584,
		54077	=>	3585,
		54078	=>	3587,
		54079	=>	3588,
		54080	=>	3590,
		54081	=>	3591,
		54082	=>	3593,
		54083	=>	3594,
		54084	=>	3595,
		54085	=>	3597,
		54086	=>	3598,
		54087	=>	3600,
		54088	=>	3601,
		54089	=>	3603,
		54090	=>	3604,
		54091	=>	3605,
		54092	=>	3607,
		54093	=>	3608,
		54094	=>	3610,
		54095	=>	3611,
		54096	=>	3613,
		54097	=>	3614,
		54098	=>	3615,
		54099	=>	3617,
		54100	=>	3618,
		54101	=>	3620,
		54102	=>	3621,
		54103	=>	3623,
		54104	=>	3624,
		54105	=>	3626,
		54106	=>	3627,
		54107	=>	3628,
		54108	=>	3630,
		54109	=>	3631,
		54110	=>	3633,
		54111	=>	3634,
		54112	=>	3636,
		54113	=>	3637,
		54114	=>	3638,
		54115	=>	3640,
		54116	=>	3641,
		54117	=>	3643,
		54118	=>	3644,
		54119	=>	3646,
		54120	=>	3647,
		54121	=>	3649,
		54122	=>	3650,
		54123	=>	3651,
		54124	=>	3653,
		54125	=>	3654,
		54126	=>	3656,
		54127	=>	3657,
		54128	=>	3659,
		54129	=>	3660,
		54130	=>	3662,
		54131	=>	3663,
		54132	=>	3664,
		54133	=>	3666,
		54134	=>	3667,
		54135	=>	3669,
		54136	=>	3670,
		54137	=>	3672,
		54138	=>	3673,
		54139	=>	3675,
		54140	=>	3676,
		54141	=>	3677,
		54142	=>	3679,
		54143	=>	3680,
		54144	=>	3682,
		54145	=>	3683,
		54146	=>	3685,
		54147	=>	3686,
		54148	=>	3688,
		54149	=>	3689,
		54150	=>	3690,
		54151	=>	3692,
		54152	=>	3693,
		54153	=>	3695,
		54154	=>	3696,
		54155	=>	3698,
		54156	=>	3699,
		54157	=>	3701,
		54158	=>	3702,
		54159	=>	3704,
		54160	=>	3705,
		54161	=>	3706,
		54162	=>	3708,
		54163	=>	3709,
		54164	=>	3711,
		54165	=>	3712,
		54166	=>	3714,
		54167	=>	3715,
		54168	=>	3717,
		54169	=>	3718,
		54170	=>	3719,
		54171	=>	3721,
		54172	=>	3722,
		54173	=>	3724,
		54174	=>	3725,
		54175	=>	3727,
		54176	=>	3728,
		54177	=>	3730,
		54178	=>	3731,
		54179	=>	3733,
		54180	=>	3734,
		54181	=>	3735,
		54182	=>	3737,
		54183	=>	3738,
		54184	=>	3740,
		54185	=>	3741,
		54186	=>	3743,
		54187	=>	3744,
		54188	=>	3746,
		54189	=>	3747,
		54190	=>	3749,
		54191	=>	3750,
		54192	=>	3752,
		54193	=>	3753,
		54194	=>	3754,
		54195	=>	3756,
		54196	=>	3757,
		54197	=>	3759,
		54198	=>	3760,
		54199	=>	3762,
		54200	=>	3763,
		54201	=>	3765,
		54202	=>	3766,
		54203	=>	3768,
		54204	=>	3769,
		54205	=>	3771,
		54206	=>	3772,
		54207	=>	3773,
		54208	=>	3775,
		54209	=>	3776,
		54210	=>	3778,
		54211	=>	3779,
		54212	=>	3781,
		54213	=>	3782,
		54214	=>	3784,
		54215	=>	3785,
		54216	=>	3787,
		54217	=>	3788,
		54218	=>	3790,
		54219	=>	3791,
		54220	=>	3792,
		54221	=>	3794,
		54222	=>	3795,
		54223	=>	3797,
		54224	=>	3798,
		54225	=>	3800,
		54226	=>	3801,
		54227	=>	3803,
		54228	=>	3804,
		54229	=>	3806,
		54230	=>	3807,
		54231	=>	3809,
		54232	=>	3810,
		54233	=>	3812,
		54234	=>	3813,
		54235	=>	3815,
		54236	=>	3816,
		54237	=>	3817,
		54238	=>	3819,
		54239	=>	3820,
		54240	=>	3822,
		54241	=>	3823,
		54242	=>	3825,
		54243	=>	3826,
		54244	=>	3828,
		54245	=>	3829,
		54246	=>	3831,
		54247	=>	3832,
		54248	=>	3834,
		54249	=>	3835,
		54250	=>	3837,
		54251	=>	3838,
		54252	=>	3840,
		54253	=>	3841,
		54254	=>	3843,
		54255	=>	3844,
		54256	=>	3845,
		54257	=>	3847,
		54258	=>	3848,
		54259	=>	3850,
		54260	=>	3851,
		54261	=>	3853,
		54262	=>	3854,
		54263	=>	3856,
		54264	=>	3857,
		54265	=>	3859,
		54266	=>	3860,
		54267	=>	3862,
		54268	=>	3863,
		54269	=>	3865,
		54270	=>	3866,
		54271	=>	3868,
		54272	=>	3869,
		54273	=>	3871,
		54274	=>	3872,
		54275	=>	3874,
		54276	=>	3875,
		54277	=>	3877,
		54278	=>	3878,
		54279	=>	3880,
		54280	=>	3881,
		54281	=>	3882,
		54282	=>	3884,
		54283	=>	3885,
		54284	=>	3887,
		54285	=>	3888,
		54286	=>	3890,
		54287	=>	3891,
		54288	=>	3893,
		54289	=>	3894,
		54290	=>	3896,
		54291	=>	3897,
		54292	=>	3899,
		54293	=>	3900,
		54294	=>	3902,
		54295	=>	3903,
		54296	=>	3905,
		54297	=>	3906,
		54298	=>	3908,
		54299	=>	3909,
		54300	=>	3911,
		54301	=>	3912,
		54302	=>	3914,
		54303	=>	3915,
		54304	=>	3917,
		54305	=>	3918,
		54306	=>	3920,
		54307	=>	3921,
		54308	=>	3923,
		54309	=>	3924,
		54310	=>	3926,
		54311	=>	3927,
		54312	=>	3929,
		54313	=>	3930,
		54314	=>	3932,
		54315	=>	3933,
		54316	=>	3935,
		54317	=>	3936,
		54318	=>	3938,
		54319	=>	3939,
		54320	=>	3941,
		54321	=>	3942,
		54322	=>	3944,
		54323	=>	3945,
		54324	=>	3947,
		54325	=>	3948,
		54326	=>	3950,
		54327	=>	3951,
		54328	=>	3952,
		54329	=>	3954,
		54330	=>	3955,
		54331	=>	3957,
		54332	=>	3958,
		54333	=>	3960,
		54334	=>	3961,
		54335	=>	3963,
		54336	=>	3964,
		54337	=>	3966,
		54338	=>	3967,
		54339	=>	3969,
		54340	=>	3970,
		54341	=>	3972,
		54342	=>	3973,
		54343	=>	3975,
		54344	=>	3976,
		54345	=>	3978,
		54346	=>	3979,
		54347	=>	3981,
		54348	=>	3982,
		54349	=>	3984,
		54350	=>	3985,
		54351	=>	3987,
		54352	=>	3988,
		54353	=>	3990,
		54354	=>	3991,
		54355	=>	3993,
		54356	=>	3994,
		54357	=>	3996,
		54358	=>	3997,
		54359	=>	3999,
		54360	=>	4000,
		54361	=>	4002,
		54362	=>	4004,
		54363	=>	4005,
		54364	=>	4007,
		54365	=>	4008,
		54366	=>	4010,
		54367	=>	4011,
		54368	=>	4013,
		54369	=>	4014,
		54370	=>	4016,
		54371	=>	4017,
		54372	=>	4019,
		54373	=>	4020,
		54374	=>	4022,
		54375	=>	4023,
		54376	=>	4025,
		54377	=>	4026,
		54378	=>	4028,
		54379	=>	4029,
		54380	=>	4031,
		54381	=>	4032,
		54382	=>	4034,
		54383	=>	4035,
		54384	=>	4037,
		54385	=>	4038,
		54386	=>	4040,
		54387	=>	4041,
		54388	=>	4043,
		54389	=>	4044,
		54390	=>	4046,
		54391	=>	4047,
		54392	=>	4049,
		54393	=>	4050,
		54394	=>	4052,
		54395	=>	4053,
		54396	=>	4055,
		54397	=>	4056,
		54398	=>	4058,
		54399	=>	4059,
		54400	=>	4061,
		54401	=>	4062,
		54402	=>	4064,
		54403	=>	4065,
		54404	=>	4067,
		54405	=>	4068,
		54406	=>	4070,
		54407	=>	4071,
		54408	=>	4073,
		54409	=>	4075,
		54410	=>	4076,
		54411	=>	4078,
		54412	=>	4079,
		54413	=>	4081,
		54414	=>	4082,
		54415	=>	4084,
		54416	=>	4085,
		54417	=>	4087,
		54418	=>	4088,
		54419	=>	4090,
		54420	=>	4091,
		54421	=>	4093,
		54422	=>	4094,
		54423	=>	4096,
		54424	=>	4097,
		54425	=>	4099,
		54426	=>	4100,
		54427	=>	4102,
		54428	=>	4103,
		54429	=>	4105,
		54430	=>	4106,
		54431	=>	4108,
		54432	=>	4109,
		54433	=>	4111,
		54434	=>	4113,
		54435	=>	4114,
		54436	=>	4116,
		54437	=>	4117,
		54438	=>	4119,
		54439	=>	4120,
		54440	=>	4122,
		54441	=>	4123,
		54442	=>	4125,
		54443	=>	4126,
		54444	=>	4128,
		54445	=>	4129,
		54446	=>	4131,
		54447	=>	4132,
		54448	=>	4134,
		54449	=>	4135,
		54450	=>	4137,
		54451	=>	4138,
		54452	=>	4140,
		54453	=>	4142,
		54454	=>	4143,
		54455	=>	4145,
		54456	=>	4146,
		54457	=>	4148,
		54458	=>	4149,
		54459	=>	4151,
		54460	=>	4152,
		54461	=>	4154,
		54462	=>	4155,
		54463	=>	4157,
		54464	=>	4158,
		54465	=>	4160,
		54466	=>	4161,
		54467	=>	4163,
		54468	=>	4164,
		54469	=>	4166,
		54470	=>	4168,
		54471	=>	4169,
		54472	=>	4171,
		54473	=>	4172,
		54474	=>	4174,
		54475	=>	4175,
		54476	=>	4177,
		54477	=>	4178,
		54478	=>	4180,
		54479	=>	4181,
		54480	=>	4183,
		54481	=>	4184,
		54482	=>	4186,
		54483	=>	4188,
		54484	=>	4189,
		54485	=>	4191,
		54486	=>	4192,
		54487	=>	4194,
		54488	=>	4195,
		54489	=>	4197,
		54490	=>	4198,
		54491	=>	4200,
		54492	=>	4201,
		54493	=>	4203,
		54494	=>	4204,
		54495	=>	4206,
		54496	=>	4208,
		54497	=>	4209,
		54498	=>	4211,
		54499	=>	4212,
		54500	=>	4214,
		54501	=>	4215,
		54502	=>	4217,
		54503	=>	4218,
		54504	=>	4220,
		54505	=>	4221,
		54506	=>	4223,
		54507	=>	4224,
		54508	=>	4226,
		54509	=>	4228,
		54510	=>	4229,
		54511	=>	4231,
		54512	=>	4232,
		54513	=>	4234,
		54514	=>	4235,
		54515	=>	4237,
		54516	=>	4238,
		54517	=>	4240,
		54518	=>	4241,
		54519	=>	4243,
		54520	=>	4245,
		54521	=>	4246,
		54522	=>	4248,
		54523	=>	4249,
		54524	=>	4251,
		54525	=>	4252,
		54526	=>	4254,
		54527	=>	4255,
		54528	=>	4257,
		54529	=>	4258,
		54530	=>	4260,
		54531	=>	4262,
		54532	=>	4263,
		54533	=>	4265,
		54534	=>	4266,
		54535	=>	4268,
		54536	=>	4269,
		54537	=>	4271,
		54538	=>	4272,
		54539	=>	4274,
		54540	=>	4276,
		54541	=>	4277,
		54542	=>	4279,
		54543	=>	4280,
		54544	=>	4282,
		54545	=>	4283,
		54546	=>	4285,
		54547	=>	4286,
		54548	=>	4288,
		54549	=>	4289,
		54550	=>	4291,
		54551	=>	4293,
		54552	=>	4294,
		54553	=>	4296,
		54554	=>	4297,
		54555	=>	4299,
		54556	=>	4300,
		54557	=>	4302,
		54558	=>	4303,
		54559	=>	4305,
		54560	=>	4307,
		54561	=>	4308,
		54562	=>	4310,
		54563	=>	4311,
		54564	=>	4313,
		54565	=>	4314,
		54566	=>	4316,
		54567	=>	4318,
		54568	=>	4319,
		54569	=>	4321,
		54570	=>	4322,
		54571	=>	4324,
		54572	=>	4325,
		54573	=>	4327,
		54574	=>	4328,
		54575	=>	4330,
		54576	=>	4332,
		54577	=>	4333,
		54578	=>	4335,
		54579	=>	4336,
		54580	=>	4338,
		54581	=>	4339,
		54582	=>	4341,
		54583	=>	4342,
		54584	=>	4344,
		54585	=>	4346,
		54586	=>	4347,
		54587	=>	4349,
		54588	=>	4350,
		54589	=>	4352,
		54590	=>	4353,
		54591	=>	4355,
		54592	=>	4357,
		54593	=>	4358,
		54594	=>	4360,
		54595	=>	4361,
		54596	=>	4363,
		54597	=>	4364,
		54598	=>	4366,
		54599	=>	4368,
		54600	=>	4369,
		54601	=>	4371,
		54602	=>	4372,
		54603	=>	4374,
		54604	=>	4375,
		54605	=>	4377,
		54606	=>	4379,
		54607	=>	4380,
		54608	=>	4382,
		54609	=>	4383,
		54610	=>	4385,
		54611	=>	4386,
		54612	=>	4388,
		54613	=>	4389,
		54614	=>	4391,
		54615	=>	4393,
		54616	=>	4394,
		54617	=>	4396,
		54618	=>	4397,
		54619	=>	4399,
		54620	=>	4400,
		54621	=>	4402,
		54622	=>	4404,
		54623	=>	4405,
		54624	=>	4407,
		54625	=>	4408,
		54626	=>	4410,
		54627	=>	4412,
		54628	=>	4413,
		54629	=>	4415,
		54630	=>	4416,
		54631	=>	4418,
		54632	=>	4419,
		54633	=>	4421,
		54634	=>	4423,
		54635	=>	4424,
		54636	=>	4426,
		54637	=>	4427,
		54638	=>	4429,
		54639	=>	4430,
		54640	=>	4432,
		54641	=>	4434,
		54642	=>	4435,
		54643	=>	4437,
		54644	=>	4438,
		54645	=>	4440,
		54646	=>	4441,
		54647	=>	4443,
		54648	=>	4445,
		54649	=>	4446,
		54650	=>	4448,
		54651	=>	4449,
		54652	=>	4451,
		54653	=>	4453,
		54654	=>	4454,
		54655	=>	4456,
		54656	=>	4457,
		54657	=>	4459,
		54658	=>	4460,
		54659	=>	4462,
		54660	=>	4464,
		54661	=>	4465,
		54662	=>	4467,
		54663	=>	4468,
		54664	=>	4470,
		54665	=>	4472,
		54666	=>	4473,
		54667	=>	4475,
		54668	=>	4476,
		54669	=>	4478,
		54670	=>	4479,
		54671	=>	4481,
		54672	=>	4483,
		54673	=>	4484,
		54674	=>	4486,
		54675	=>	4487,
		54676	=>	4489,
		54677	=>	4491,
		54678	=>	4492,
		54679	=>	4494,
		54680	=>	4495,
		54681	=>	4497,
		54682	=>	4498,
		54683	=>	4500,
		54684	=>	4502,
		54685	=>	4503,
		54686	=>	4505,
		54687	=>	4506,
		54688	=>	4508,
		54689	=>	4510,
		54690	=>	4511,
		54691	=>	4513,
		54692	=>	4514,
		54693	=>	4516,
		54694	=>	4518,
		54695	=>	4519,
		54696	=>	4521,
		54697	=>	4522,
		54698	=>	4524,
		54699	=>	4526,
		54700	=>	4527,
		54701	=>	4529,
		54702	=>	4530,
		54703	=>	4532,
		54704	=>	4533,
		54705	=>	4535,
		54706	=>	4537,
		54707	=>	4538,
		54708	=>	4540,
		54709	=>	4541,
		54710	=>	4543,
		54711	=>	4545,
		54712	=>	4546,
		54713	=>	4548,
		54714	=>	4549,
		54715	=>	4551,
		54716	=>	4553,
		54717	=>	4554,
		54718	=>	4556,
		54719	=>	4557,
		54720	=>	4559,
		54721	=>	4561,
		54722	=>	4562,
		54723	=>	4564,
		54724	=>	4565,
		54725	=>	4567,
		54726	=>	4569,
		54727	=>	4570,
		54728	=>	4572,
		54729	=>	4573,
		54730	=>	4575,
		54731	=>	4577,
		54732	=>	4578,
		54733	=>	4580,
		54734	=>	4581,
		54735	=>	4583,
		54736	=>	4585,
		54737	=>	4586,
		54738	=>	4588,
		54739	=>	4589,
		54740	=>	4591,
		54741	=>	4593,
		54742	=>	4594,
		54743	=>	4596,
		54744	=>	4597,
		54745	=>	4599,
		54746	=>	4601,
		54747	=>	4602,
		54748	=>	4604,
		54749	=>	4606,
		54750	=>	4607,
		54751	=>	4609,
		54752	=>	4610,
		54753	=>	4612,
		54754	=>	4614,
		54755	=>	4615,
		54756	=>	4617,
		54757	=>	4618,
		54758	=>	4620,
		54759	=>	4622,
		54760	=>	4623,
		54761	=>	4625,
		54762	=>	4626,
		54763	=>	4628,
		54764	=>	4630,
		54765	=>	4631,
		54766	=>	4633,
		54767	=>	4634,
		54768	=>	4636,
		54769	=>	4638,
		54770	=>	4639,
		54771	=>	4641,
		54772	=>	4643,
		54773	=>	4644,
		54774	=>	4646,
		54775	=>	4647,
		54776	=>	4649,
		54777	=>	4651,
		54778	=>	4652,
		54779	=>	4654,
		54780	=>	4655,
		54781	=>	4657,
		54782	=>	4659,
		54783	=>	4660,
		54784	=>	4662,
		54785	=>	4663,
		54786	=>	4665,
		54787	=>	4667,
		54788	=>	4668,
		54789	=>	4670,
		54790	=>	4672,
		54791	=>	4673,
		54792	=>	4675,
		54793	=>	4676,
		54794	=>	4678,
		54795	=>	4680,
		54796	=>	4681,
		54797	=>	4683,
		54798	=>	4685,
		54799	=>	4686,
		54800	=>	4688,
		54801	=>	4689,
		54802	=>	4691,
		54803	=>	4693,
		54804	=>	4694,
		54805	=>	4696,
		54806	=>	4697,
		54807	=>	4699,
		54808	=>	4701,
		54809	=>	4702,
		54810	=>	4704,
		54811	=>	4706,
		54812	=>	4707,
		54813	=>	4709,
		54814	=>	4710,
		54815	=>	4712,
		54816	=>	4714,
		54817	=>	4715,
		54818	=>	4717,
		54819	=>	4719,
		54820	=>	4720,
		54821	=>	4722,
		54822	=>	4723,
		54823	=>	4725,
		54824	=>	4727,
		54825	=>	4728,
		54826	=>	4730,
		54827	=>	4732,
		54828	=>	4733,
		54829	=>	4735,
		54830	=>	4736,
		54831	=>	4738,
		54832	=>	4740,
		54833	=>	4741,
		54834	=>	4743,
		54835	=>	4745,
		54836	=>	4746,
		54837	=>	4748,
		54838	=>	4749,
		54839	=>	4751,
		54840	=>	4753,
		54841	=>	4754,
		54842	=>	4756,
		54843	=>	4758,
		54844	=>	4759,
		54845	=>	4761,
		54846	=>	4763,
		54847	=>	4764,
		54848	=>	4766,
		54849	=>	4767,
		54850	=>	4769,
		54851	=>	4771,
		54852	=>	4772,
		54853	=>	4774,
		54854	=>	4776,
		54855	=>	4777,
		54856	=>	4779,
		54857	=>	4780,
		54858	=>	4782,
		54859	=>	4784,
		54860	=>	4785,
		54861	=>	4787,
		54862	=>	4789,
		54863	=>	4790,
		54864	=>	4792,
		54865	=>	4794,
		54866	=>	4795,
		54867	=>	4797,
		54868	=>	4798,
		54869	=>	4800,
		54870	=>	4802,
		54871	=>	4803,
		54872	=>	4805,
		54873	=>	4807,
		54874	=>	4808,
		54875	=>	4810,
		54876	=>	4812,
		54877	=>	4813,
		54878	=>	4815,
		54879	=>	4816,
		54880	=>	4818,
		54881	=>	4820,
		54882	=>	4821,
		54883	=>	4823,
		54884	=>	4825,
		54885	=>	4826,
		54886	=>	4828,
		54887	=>	4830,
		54888	=>	4831,
		54889	=>	4833,
		54890	=>	4835,
		54891	=>	4836,
		54892	=>	4838,
		54893	=>	4839,
		54894	=>	4841,
		54895	=>	4843,
		54896	=>	4844,
		54897	=>	4846,
		54898	=>	4848,
		54899	=>	4849,
		54900	=>	4851,
		54901	=>	4853,
		54902	=>	4854,
		54903	=>	4856,
		54904	=>	4858,
		54905	=>	4859,
		54906	=>	4861,
		54907	=>	4862,
		54908	=>	4864,
		54909	=>	4866,
		54910	=>	4867,
		54911	=>	4869,
		54912	=>	4871,
		54913	=>	4872,
		54914	=>	4874,
		54915	=>	4876,
		54916	=>	4877,
		54917	=>	4879,
		54918	=>	4881,
		54919	=>	4882,
		54920	=>	4884,
		54921	=>	4886,
		54922	=>	4887,
		54923	=>	4889,
		54924	=>	4891,
		54925	=>	4892,
		54926	=>	4894,
		54927	=>	4895,
		54928	=>	4897,
		54929	=>	4899,
		54930	=>	4900,
		54931	=>	4902,
		54932	=>	4904,
		54933	=>	4905,
		54934	=>	4907,
		54935	=>	4909,
		54936	=>	4910,
		54937	=>	4912,
		54938	=>	4914,
		54939	=>	4915,
		54940	=>	4917,
		54941	=>	4919,
		54942	=>	4920,
		54943	=>	4922,
		54944	=>	4924,
		54945	=>	4925,
		54946	=>	4927,
		54947	=>	4929,
		54948	=>	4930,
		54949	=>	4932,
		54950	=>	4934,
		54951	=>	4935,
		54952	=>	4937,
		54953	=>	4939,
		54954	=>	4940,
		54955	=>	4942,
		54956	=>	4943,
		54957	=>	4945,
		54958	=>	4947,
		54959	=>	4948,
		54960	=>	4950,
		54961	=>	4952,
		54962	=>	4953,
		54963	=>	4955,
		54964	=>	4957,
		54965	=>	4958,
		54966	=>	4960,
		54967	=>	4962,
		54968	=>	4963,
		54969	=>	4965,
		54970	=>	4967,
		54971	=>	4968,
		54972	=>	4970,
		54973	=>	4972,
		54974	=>	4973,
		54975	=>	4975,
		54976	=>	4977,
		54977	=>	4978,
		54978	=>	4980,
		54979	=>	4982,
		54980	=>	4983,
		54981	=>	4985,
		54982	=>	4987,
		54983	=>	4988,
		54984	=>	4990,
		54985	=>	4992,
		54986	=>	4993,
		54987	=>	4995,
		54988	=>	4997,
		54989	=>	4998,
		54990	=>	5000,
		54991	=>	5002,
		54992	=>	5003,
		54993	=>	5005,
		54994	=>	5007,
		54995	=>	5008,
		54996	=>	5010,
		54997	=>	5012,
		54998	=>	5013,
		54999	=>	5015,
		55000	=>	5017,
		55001	=>	5018,
		55002	=>	5020,
		55003	=>	5022,
		55004	=>	5023,
		55005	=>	5025,
		55006	=>	5027,
		55007	=>	5028,
		55008	=>	5030,
		55009	=>	5032,
		55010	=>	5033,
		55011	=>	5035,
		55012	=>	5037,
		55013	=>	5038,
		55014	=>	5040,
		55015	=>	5042,
		55016	=>	5043,
		55017	=>	5045,
		55018	=>	5047,
		55019	=>	5049,
		55020	=>	5050,
		55021	=>	5052,
		55022	=>	5054,
		55023	=>	5055,
		55024	=>	5057,
		55025	=>	5059,
		55026	=>	5060,
		55027	=>	5062,
		55028	=>	5064,
		55029	=>	5065,
		55030	=>	5067,
		55031	=>	5069,
		55032	=>	5070,
		55033	=>	5072,
		55034	=>	5074,
		55035	=>	5075,
		55036	=>	5077,
		55037	=>	5079,
		55038	=>	5080,
		55039	=>	5082,
		55040	=>	5084,
		55041	=>	5085,
		55042	=>	5087,
		55043	=>	5089,
		55044	=>	5090,
		55045	=>	5092,
		55046	=>	5094,
		55047	=>	5096,
		55048	=>	5097,
		55049	=>	5099,
		55050	=>	5101,
		55051	=>	5102,
		55052	=>	5104,
		55053	=>	5106,
		55054	=>	5107,
		55055	=>	5109,
		55056	=>	5111,
		55057	=>	5112,
		55058	=>	5114,
		55059	=>	5116,
		55060	=>	5117,
		55061	=>	5119,
		55062	=>	5121,
		55063	=>	5122,
		55064	=>	5124,
		55065	=>	5126,
		55066	=>	5128,
		55067	=>	5129,
		55068	=>	5131,
		55069	=>	5133,
		55070	=>	5134,
		55071	=>	5136,
		55072	=>	5138,
		55073	=>	5139,
		55074	=>	5141,
		55075	=>	5143,
		55076	=>	5144,
		55077	=>	5146,
		55078	=>	5148,
		55079	=>	5150,
		55080	=>	5151,
		55081	=>	5153,
		55082	=>	5155,
		55083	=>	5156,
		55084	=>	5158,
		55085	=>	5160,
		55086	=>	5161,
		55087	=>	5163,
		55088	=>	5165,
		55089	=>	5166,
		55090	=>	5168,
		55091	=>	5170,
		55092	=>	5172,
		55093	=>	5173,
		55094	=>	5175,
		55095	=>	5177,
		55096	=>	5178,
		55097	=>	5180,
		55098	=>	5182,
		55099	=>	5183,
		55100	=>	5185,
		55101	=>	5187,
		55102	=>	5188,
		55103	=>	5190,
		55104	=>	5192,
		55105	=>	5194,
		55106	=>	5195,
		55107	=>	5197,
		55108	=>	5199,
		55109	=>	5200,
		55110	=>	5202,
		55111	=>	5204,
		55112	=>	5205,
		55113	=>	5207,
		55114	=>	5209,
		55115	=>	5211,
		55116	=>	5212,
		55117	=>	5214,
		55118	=>	5216,
		55119	=>	5217,
		55120	=>	5219,
		55121	=>	5221,
		55122	=>	5222,
		55123	=>	5224,
		55124	=>	5226,
		55125	=>	5228,
		55126	=>	5229,
		55127	=>	5231,
		55128	=>	5233,
		55129	=>	5234,
		55130	=>	5236,
		55131	=>	5238,
		55132	=>	5239,
		55133	=>	5241,
		55134	=>	5243,
		55135	=>	5245,
		55136	=>	5246,
		55137	=>	5248,
		55138	=>	5250,
		55139	=>	5251,
		55140	=>	5253,
		55141	=>	5255,
		55142	=>	5257,
		55143	=>	5258,
		55144	=>	5260,
		55145	=>	5262,
		55146	=>	5263,
		55147	=>	5265,
		55148	=>	5267,
		55149	=>	5268,
		55150	=>	5270,
		55151	=>	5272,
		55152	=>	5274,
		55153	=>	5275,
		55154	=>	5277,
		55155	=>	5279,
		55156	=>	5280,
		55157	=>	5282,
		55158	=>	5284,
		55159	=>	5286,
		55160	=>	5287,
		55161	=>	5289,
		55162	=>	5291,
		55163	=>	5292,
		55164	=>	5294,
		55165	=>	5296,
		55166	=>	5298,
		55167	=>	5299,
		55168	=>	5301,
		55169	=>	5303,
		55170	=>	5304,
		55171	=>	5306,
		55172	=>	5308,
		55173	=>	5310,
		55174	=>	5311,
		55175	=>	5313,
		55176	=>	5315,
		55177	=>	5316,
		55178	=>	5318,
		55179	=>	5320,
		55180	=>	5322,
		55181	=>	5323,
		55182	=>	5325,
		55183	=>	5327,
		55184	=>	5328,
		55185	=>	5330,
		55186	=>	5332,
		55187	=>	5334,
		55188	=>	5335,
		55189	=>	5337,
		55190	=>	5339,
		55191	=>	5340,
		55192	=>	5342,
		55193	=>	5344,
		55194	=>	5346,
		55195	=>	5347,
		55196	=>	5349,
		55197	=>	5351,
		55198	=>	5352,
		55199	=>	5354,
		55200	=>	5356,
		55201	=>	5358,
		55202	=>	5359,
		55203	=>	5361,
		55204	=>	5363,
		55205	=>	5365,
		55206	=>	5366,
		55207	=>	5368,
		55208	=>	5370,
		55209	=>	5371,
		55210	=>	5373,
		55211	=>	5375,
		55212	=>	5377,
		55213	=>	5378,
		55214	=>	5380,
		55215	=>	5382,
		55216	=>	5383,
		55217	=>	5385,
		55218	=>	5387,
		55219	=>	5389,
		55220	=>	5390,
		55221	=>	5392,
		55222	=>	5394,
		55223	=>	5396,
		55224	=>	5397,
		55225	=>	5399,
		55226	=>	5401,
		55227	=>	5402,
		55228	=>	5404,
		55229	=>	5406,
		55230	=>	5408,
		55231	=>	5409,
		55232	=>	5411,
		55233	=>	5413,
		55234	=>	5415,
		55235	=>	5416,
		55236	=>	5418,
		55237	=>	5420,
		55238	=>	5422,
		55239	=>	5423,
		55240	=>	5425,
		55241	=>	5427,
		55242	=>	5428,
		55243	=>	5430,
		55244	=>	5432,
		55245	=>	5434,
		55246	=>	5435,
		55247	=>	5437,
		55248	=>	5439,
		55249	=>	5441,
		55250	=>	5442,
		55251	=>	5444,
		55252	=>	5446,
		55253	=>	5448,
		55254	=>	5449,
		55255	=>	5451,
		55256	=>	5453,
		55257	=>	5454,
		55258	=>	5456,
		55259	=>	5458,
		55260	=>	5460,
		55261	=>	5461,
		55262	=>	5463,
		55263	=>	5465,
		55264	=>	5467,
		55265	=>	5468,
		55266	=>	5470,
		55267	=>	5472,
		55268	=>	5474,
		55269	=>	5475,
		55270	=>	5477,
		55271	=>	5479,
		55272	=>	5481,
		55273	=>	5482,
		55274	=>	5484,
		55275	=>	5486,
		55276	=>	5487,
		55277	=>	5489,
		55278	=>	5491,
		55279	=>	5493,
		55280	=>	5494,
		55281	=>	5496,
		55282	=>	5498,
		55283	=>	5500,
		55284	=>	5501,
		55285	=>	5503,
		55286	=>	5505,
		55287	=>	5507,
		55288	=>	5508,
		55289	=>	5510,
		55290	=>	5512,
		55291	=>	5514,
		55292	=>	5515,
		55293	=>	5517,
		55294	=>	5519,
		55295	=>	5521,
		55296	=>	5522,
		55297	=>	5524,
		55298	=>	5526,
		55299	=>	5528,
		55300	=>	5529,
		55301	=>	5531,
		55302	=>	5533,
		55303	=>	5535,
		55304	=>	5536,
		55305	=>	5538,
		55306	=>	5540,
		55307	=>	5542,
		55308	=>	5543,
		55309	=>	5545,
		55310	=>	5547,
		55311	=>	5549,
		55312	=>	5550,
		55313	=>	5552,
		55314	=>	5554,
		55315	=>	5556,
		55316	=>	5557,
		55317	=>	5559,
		55318	=>	5561,
		55319	=>	5563,
		55320	=>	5564,
		55321	=>	5566,
		55322	=>	5568,
		55323	=>	5570,
		55324	=>	5571,
		55325	=>	5573,
		55326	=>	5575,
		55327	=>	5577,
		55328	=>	5578,
		55329	=>	5580,
		55330	=>	5582,
		55331	=>	5584,
		55332	=>	5585,
		55333	=>	5587,
		55334	=>	5589,
		55335	=>	5591,
		55336	=>	5592,
		55337	=>	5594,
		55338	=>	5596,
		55339	=>	5598,
		55340	=>	5599,
		55341	=>	5601,
		55342	=>	5603,
		55343	=>	5605,
		55344	=>	5606,
		55345	=>	5608,
		55346	=>	5610,
		55347	=>	5612,
		55348	=>	5613,
		55349	=>	5615,
		55350	=>	5617,
		55351	=>	5619,
		55352	=>	5620,
		55353	=>	5622,
		55354	=>	5624,
		55355	=>	5626,
		55356	=>	5627,
		55357	=>	5629,
		55358	=>	5631,
		55359	=>	5633,
		55360	=>	5635,
		55361	=>	5636,
		55362	=>	5638,
		55363	=>	5640,
		55364	=>	5642,
		55365	=>	5643,
		55366	=>	5645,
		55367	=>	5647,
		55368	=>	5649,
		55369	=>	5650,
		55370	=>	5652,
		55371	=>	5654,
		55372	=>	5656,
		55373	=>	5657,
		55374	=>	5659,
		55375	=>	5661,
		55376	=>	5663,
		55377	=>	5665,
		55378	=>	5666,
		55379	=>	5668,
		55380	=>	5670,
		55381	=>	5672,
		55382	=>	5673,
		55383	=>	5675,
		55384	=>	5677,
		55385	=>	5679,
		55386	=>	5680,
		55387	=>	5682,
		55388	=>	5684,
		55389	=>	5686,
		55390	=>	5687,
		55391	=>	5689,
		55392	=>	5691,
		55393	=>	5693,
		55394	=>	5695,
		55395	=>	5696,
		55396	=>	5698,
		55397	=>	5700,
		55398	=>	5702,
		55399	=>	5703,
		55400	=>	5705,
		55401	=>	5707,
		55402	=>	5709,
		55403	=>	5711,
		55404	=>	5712,
		55405	=>	5714,
		55406	=>	5716,
		55407	=>	5718,
		55408	=>	5719,
		55409	=>	5721,
		55410	=>	5723,
		55411	=>	5725,
		55412	=>	5726,
		55413	=>	5728,
		55414	=>	5730,
		55415	=>	5732,
		55416	=>	5734,
		55417	=>	5735,
		55418	=>	5737,
		55419	=>	5739,
		55420	=>	5741,
		55421	=>	5742,
		55422	=>	5744,
		55423	=>	5746,
		55424	=>	5748,
		55425	=>	5750,
		55426	=>	5751,
		55427	=>	5753,
		55428	=>	5755,
		55429	=>	5757,
		55430	=>	5758,
		55431	=>	5760,
		55432	=>	5762,
		55433	=>	5764,
		55434	=>	5766,
		55435	=>	5767,
		55436	=>	5769,
		55437	=>	5771,
		55438	=>	5773,
		55439	=>	5774,
		55440	=>	5776,
		55441	=>	5778,
		55442	=>	5780,
		55443	=>	5782,
		55444	=>	5783,
		55445	=>	5785,
		55446	=>	5787,
		55447	=>	5789,
		55448	=>	5790,
		55449	=>	5792,
		55450	=>	5794,
		55451	=>	5796,
		55452	=>	5798,
		55453	=>	5799,
		55454	=>	5801,
		55455	=>	5803,
		55456	=>	5805,
		55457	=>	5807,
		55458	=>	5808,
		55459	=>	5810,
		55460	=>	5812,
		55461	=>	5814,
		55462	=>	5815,
		55463	=>	5817,
		55464	=>	5819,
		55465	=>	5821,
		55466	=>	5823,
		55467	=>	5824,
		55468	=>	5826,
		55469	=>	5828,
		55470	=>	5830,
		55471	=>	5832,
		55472	=>	5833,
		55473	=>	5835,
		55474	=>	5837,
		55475	=>	5839,
		55476	=>	5841,
		55477	=>	5842,
		55478	=>	5844,
		55479	=>	5846,
		55480	=>	5848,
		55481	=>	5849,
		55482	=>	5851,
		55483	=>	5853,
		55484	=>	5855,
		55485	=>	5857,
		55486	=>	5858,
		55487	=>	5860,
		55488	=>	5862,
		55489	=>	5864,
		55490	=>	5866,
		55491	=>	5867,
		55492	=>	5869,
		55493	=>	5871,
		55494	=>	5873,
		55495	=>	5875,
		55496	=>	5876,
		55497	=>	5878,
		55498	=>	5880,
		55499	=>	5882,
		55500	=>	5884,
		55501	=>	5885,
		55502	=>	5887,
		55503	=>	5889,
		55504	=>	5891,
		55505	=>	5893,
		55506	=>	5894,
		55507	=>	5896,
		55508	=>	5898,
		55509	=>	5900,
		55510	=>	5902,
		55511	=>	5903,
		55512	=>	5905,
		55513	=>	5907,
		55514	=>	5909,
		55515	=>	5911,
		55516	=>	5912,
		55517	=>	5914,
		55518	=>	5916,
		55519	=>	5918,
		55520	=>	5920,
		55521	=>	5921,
		55522	=>	5923,
		55523	=>	5925,
		55524	=>	5927,
		55525	=>	5929,
		55526	=>	5930,
		55527	=>	5932,
		55528	=>	5934,
		55529	=>	5936,
		55530	=>	5938,
		55531	=>	5939,
		55532	=>	5941,
		55533	=>	5943,
		55534	=>	5945,
		55535	=>	5947,
		55536	=>	5948,
		55537	=>	5950,
		55538	=>	5952,
		55539	=>	5954,
		55540	=>	5956,
		55541	=>	5957,
		55542	=>	5959,
		55543	=>	5961,
		55544	=>	5963,
		55545	=>	5965,
		55546	=>	5966,
		55547	=>	5968,
		55548	=>	5970,
		55549	=>	5972,
		55550	=>	5974,
		55551	=>	5975,
		55552	=>	5977,
		55553	=>	5979,
		55554	=>	5981,
		55555	=>	5983,
		55556	=>	5985,
		55557	=>	5986,
		55558	=>	5988,
		55559	=>	5990,
		55560	=>	5992,
		55561	=>	5994,
		55562	=>	5995,
		55563	=>	5997,
		55564	=>	5999,
		55565	=>	6001,
		55566	=>	6003,
		55567	=>	6004,
		55568	=>	6006,
		55569	=>	6008,
		55570	=>	6010,
		55571	=>	6012,
		55572	=>	6014,
		55573	=>	6015,
		55574	=>	6017,
		55575	=>	6019,
		55576	=>	6021,
		55577	=>	6023,
		55578	=>	6024,
		55579	=>	6026,
		55580	=>	6028,
		55581	=>	6030,
		55582	=>	6032,
		55583	=>	6033,
		55584	=>	6035,
		55585	=>	6037,
		55586	=>	6039,
		55587	=>	6041,
		55588	=>	6043,
		55589	=>	6044,
		55590	=>	6046,
		55591	=>	6048,
		55592	=>	6050,
		55593	=>	6052,
		55594	=>	6053,
		55595	=>	6055,
		55596	=>	6057,
		55597	=>	6059,
		55598	=>	6061,
		55599	=>	6063,
		55600	=>	6064,
		55601	=>	6066,
		55602	=>	6068,
		55603	=>	6070,
		55604	=>	6072,
		55605	=>	6074,
		55606	=>	6075,
		55607	=>	6077,
		55608	=>	6079,
		55609	=>	6081,
		55610	=>	6083,
		55611	=>	6084,
		55612	=>	6086,
		55613	=>	6088,
		55614	=>	6090,
		55615	=>	6092,
		55616	=>	6094,
		55617	=>	6095,
		55618	=>	6097,
		55619	=>	6099,
		55620	=>	6101,
		55621	=>	6103,
		55622	=>	6105,
		55623	=>	6106,
		55624	=>	6108,
		55625	=>	6110,
		55626	=>	6112,
		55627	=>	6114,
		55628	=>	6115,
		55629	=>	6117,
		55630	=>	6119,
		55631	=>	6121,
		55632	=>	6123,
		55633	=>	6125,
		55634	=>	6126,
		55635	=>	6128,
		55636	=>	6130,
		55637	=>	6132,
		55638	=>	6134,
		55639	=>	6136,
		55640	=>	6137,
		55641	=>	6139,
		55642	=>	6141,
		55643	=>	6143,
		55644	=>	6145,
		55645	=>	6147,
		55646	=>	6148,
		55647	=>	6150,
		55648	=>	6152,
		55649	=>	6154,
		55650	=>	6156,
		55651	=>	6158,
		55652	=>	6159,
		55653	=>	6161,
		55654	=>	6163,
		55655	=>	6165,
		55656	=>	6167,
		55657	=>	6169,
		55658	=>	6170,
		55659	=>	6172,
		55660	=>	6174,
		55661	=>	6176,
		55662	=>	6178,
		55663	=>	6180,
		55664	=>	6181,
		55665	=>	6183,
		55666	=>	6185,
		55667	=>	6187,
		55668	=>	6189,
		55669	=>	6191,
		55670	=>	6192,
		55671	=>	6194,
		55672	=>	6196,
		55673	=>	6198,
		55674	=>	6200,
		55675	=>	6202,
		55676	=>	6203,
		55677	=>	6205,
		55678	=>	6207,
		55679	=>	6209,
		55680	=>	6211,
		55681	=>	6213,
		55682	=>	6215,
		55683	=>	6216,
		55684	=>	6218,
		55685	=>	6220,
		55686	=>	6222,
		55687	=>	6224,
		55688	=>	6226,
		55689	=>	6227,
		55690	=>	6229,
		55691	=>	6231,
		55692	=>	6233,
		55693	=>	6235,
		55694	=>	6237,
		55695	=>	6238,
		55696	=>	6240,
		55697	=>	6242,
		55698	=>	6244,
		55699	=>	6246,
		55700	=>	6248,
		55701	=>	6250,
		55702	=>	6251,
		55703	=>	6253,
		55704	=>	6255,
		55705	=>	6257,
		55706	=>	6259,
		55707	=>	6261,
		55708	=>	6262,
		55709	=>	6264,
		55710	=>	6266,
		55711	=>	6268,
		55712	=>	6270,
		55713	=>	6272,
		55714	=>	6274,
		55715	=>	6275,
		55716	=>	6277,
		55717	=>	6279,
		55718	=>	6281,
		55719	=>	6283,
		55720	=>	6285,
		55721	=>	6287,
		55722	=>	6288,
		55723	=>	6290,
		55724	=>	6292,
		55725	=>	6294,
		55726	=>	6296,
		55727	=>	6298,
		55728	=>	6299,
		55729	=>	6301,
		55730	=>	6303,
		55731	=>	6305,
		55732	=>	6307,
		55733	=>	6309,
		55734	=>	6311,
		55735	=>	6312,
		55736	=>	6314,
		55737	=>	6316,
		55738	=>	6318,
		55739	=>	6320,
		55740	=>	6322,
		55741	=>	6324,
		55742	=>	6325,
		55743	=>	6327,
		55744	=>	6329,
		55745	=>	6331,
		55746	=>	6333,
		55747	=>	6335,
		55748	=>	6337,
		55749	=>	6338,
		55750	=>	6340,
		55751	=>	6342,
		55752	=>	6344,
		55753	=>	6346,
		55754	=>	6348,
		55755	=>	6350,
		55756	=>	6351,
		55757	=>	6353,
		55758	=>	6355,
		55759	=>	6357,
		55760	=>	6359,
		55761	=>	6361,
		55762	=>	6363,
		55763	=>	6364,
		55764	=>	6366,
		55765	=>	6368,
		55766	=>	6370,
		55767	=>	6372,
		55768	=>	6374,
		55769	=>	6376,
		55770	=>	6377,
		55771	=>	6379,
		55772	=>	6381,
		55773	=>	6383,
		55774	=>	6385,
		55775	=>	6387,
		55776	=>	6389,
		55777	=>	6390,
		55778	=>	6392,
		55779	=>	6394,
		55780	=>	6396,
		55781	=>	6398,
		55782	=>	6400,
		55783	=>	6402,
		55784	=>	6404,
		55785	=>	6405,
		55786	=>	6407,
		55787	=>	6409,
		55788	=>	6411,
		55789	=>	6413,
		55790	=>	6415,
		55791	=>	6417,
		55792	=>	6418,
		55793	=>	6420,
		55794	=>	6422,
		55795	=>	6424,
		55796	=>	6426,
		55797	=>	6428,
		55798	=>	6430,
		55799	=>	6432,
		55800	=>	6433,
		55801	=>	6435,
		55802	=>	6437,
		55803	=>	6439,
		55804	=>	6441,
		55805	=>	6443,
		55806	=>	6445,
		55807	=>	6447,
		55808	=>	6448,
		55809	=>	6450,
		55810	=>	6452,
		55811	=>	6454,
		55812	=>	6456,
		55813	=>	6458,
		55814	=>	6460,
		55815	=>	6462,
		55816	=>	6463,
		55817	=>	6465,
		55818	=>	6467,
		55819	=>	6469,
		55820	=>	6471,
		55821	=>	6473,
		55822	=>	6475,
		55823	=>	6476,
		55824	=>	6478,
		55825	=>	6480,
		55826	=>	6482,
		55827	=>	6484,
		55828	=>	6486,
		55829	=>	6488,
		55830	=>	6490,
		55831	=>	6492,
		55832	=>	6493,
		55833	=>	6495,
		55834	=>	6497,
		55835	=>	6499,
		55836	=>	6501,
		55837	=>	6503,
		55838	=>	6505,
		55839	=>	6507,
		55840	=>	6508,
		55841	=>	6510,
		55842	=>	6512,
		55843	=>	6514,
		55844	=>	6516,
		55845	=>	6518,
		55846	=>	6520,
		55847	=>	6522,
		55848	=>	6523,
		55849	=>	6525,
		55850	=>	6527,
		55851	=>	6529,
		55852	=>	6531,
		55853	=>	6533,
		55854	=>	6535,
		55855	=>	6537,
		55856	=>	6539,
		55857	=>	6540,
		55858	=>	6542,
		55859	=>	6544,
		55860	=>	6546,
		55861	=>	6548,
		55862	=>	6550,
		55863	=>	6552,
		55864	=>	6554,
		55865	=>	6555,
		55866	=>	6557,
		55867	=>	6559,
		55868	=>	6561,
		55869	=>	6563,
		55870	=>	6565,
		55871	=>	6567,
		55872	=>	6569,
		55873	=>	6571,
		55874	=>	6572,
		55875	=>	6574,
		55876	=>	6576,
		55877	=>	6578,
		55878	=>	6580,
		55879	=>	6582,
		55880	=>	6584,
		55881	=>	6586,
		55882	=>	6588,
		55883	=>	6589,
		55884	=>	6591,
		55885	=>	6593,
		55886	=>	6595,
		55887	=>	6597,
		55888	=>	6599,
		55889	=>	6601,
		55890	=>	6603,
		55891	=>	6605,
		55892	=>	6606,
		55893	=>	6608,
		55894	=>	6610,
		55895	=>	6612,
		55896	=>	6614,
		55897	=>	6616,
		55898	=>	6618,
		55899	=>	6620,
		55900	=>	6622,
		55901	=>	6623,
		55902	=>	6625,
		55903	=>	6627,
		55904	=>	6629,
		55905	=>	6631,
		55906	=>	6633,
		55907	=>	6635,
		55908	=>	6637,
		55909	=>	6639,
		55910	=>	6641,
		55911	=>	6642,
		55912	=>	6644,
		55913	=>	6646,
		55914	=>	6648,
		55915	=>	6650,
		55916	=>	6652,
		55917	=>	6654,
		55918	=>	6656,
		55919	=>	6658,
		55920	=>	6660,
		55921	=>	6661,
		55922	=>	6663,
		55923	=>	6665,
		55924	=>	6667,
		55925	=>	6669,
		55926	=>	6671,
		55927	=>	6673,
		55928	=>	6675,
		55929	=>	6677,
		55930	=>	6679,
		55931	=>	6680,
		55932	=>	6682,
		55933	=>	6684,
		55934	=>	6686,
		55935	=>	6688,
		55936	=>	6690,
		55937	=>	6692,
		55938	=>	6694,
		55939	=>	6696,
		55940	=>	6698,
		55941	=>	6699,
		55942	=>	6701,
		55943	=>	6703,
		55944	=>	6705,
		55945	=>	6707,
		55946	=>	6709,
		55947	=>	6711,
		55948	=>	6713,
		55949	=>	6715,
		55950	=>	6717,
		55951	=>	6718,
		55952	=>	6720,
		55953	=>	6722,
		55954	=>	6724,
		55955	=>	6726,
		55956	=>	6728,
		55957	=>	6730,
		55958	=>	6732,
		55959	=>	6734,
		55960	=>	6736,
		55961	=>	6738,
		55962	=>	6739,
		55963	=>	6741,
		55964	=>	6743,
		55965	=>	6745,
		55966	=>	6747,
		55967	=>	6749,
		55968	=>	6751,
		55969	=>	6753,
		55970	=>	6755,
		55971	=>	6757,
		55972	=>	6759,
		55973	=>	6760,
		55974	=>	6762,
		55975	=>	6764,
		55976	=>	6766,
		55977	=>	6768,
		55978	=>	6770,
		55979	=>	6772,
		55980	=>	6774,
		55981	=>	6776,
		55982	=>	6778,
		55983	=>	6780,
		55984	=>	6781,
		55985	=>	6783,
		55986	=>	6785,
		55987	=>	6787,
		55988	=>	6789,
		55989	=>	6791,
		55990	=>	6793,
		55991	=>	6795,
		55992	=>	6797,
		55993	=>	6799,
		55994	=>	6801,
		55995	=>	6803,
		55996	=>	6804,
		55997	=>	6806,
		55998	=>	6808,
		55999	=>	6810,
		56000	=>	6812,
		56001	=>	6814,
		56002	=>	6816,
		56003	=>	6818,
		56004	=>	6820,
		56005	=>	6822,
		56006	=>	6824,
		56007	=>	6826,
		56008	=>	6827,
		56009	=>	6829,
		56010	=>	6831,
		56011	=>	6833,
		56012	=>	6835,
		56013	=>	6837,
		56014	=>	6839,
		56015	=>	6841,
		56016	=>	6843,
		56017	=>	6845,
		56018	=>	6847,
		56019	=>	6849,
		56020	=>	6851,
		56021	=>	6852,
		56022	=>	6854,
		56023	=>	6856,
		56024	=>	6858,
		56025	=>	6860,
		56026	=>	6862,
		56027	=>	6864,
		56028	=>	6866,
		56029	=>	6868,
		56030	=>	6870,
		56031	=>	6872,
		56032	=>	6874,
		56033	=>	6876,
		56034	=>	6877,
		56035	=>	6879,
		56036	=>	6881,
		56037	=>	6883,
		56038	=>	6885,
		56039	=>	6887,
		56040	=>	6889,
		56041	=>	6891,
		56042	=>	6893,
		56043	=>	6895,
		56044	=>	6897,
		56045	=>	6899,
		56046	=>	6901,
		56047	=>	6903,
		56048	=>	6904,
		56049	=>	6906,
		56050	=>	6908,
		56051	=>	6910,
		56052	=>	6912,
		56053	=>	6914,
		56054	=>	6916,
		56055	=>	6918,
		56056	=>	6920,
		56057	=>	6922,
		56058	=>	6924,
		56059	=>	6926,
		56060	=>	6928,
		56061	=>	6930,
		56062	=>	6931,
		56063	=>	6933,
		56064	=>	6935,
		56065	=>	6937,
		56066	=>	6939,
		56067	=>	6941,
		56068	=>	6943,
		56069	=>	6945,
		56070	=>	6947,
		56071	=>	6949,
		56072	=>	6951,
		56073	=>	6953,
		56074	=>	6955,
		56075	=>	6957,
		56076	=>	6959,
		56077	=>	6961,
		56078	=>	6962,
		56079	=>	6964,
		56080	=>	6966,
		56081	=>	6968,
		56082	=>	6970,
		56083	=>	6972,
		56084	=>	6974,
		56085	=>	6976,
		56086	=>	6978,
		56087	=>	6980,
		56088	=>	6982,
		56089	=>	6984,
		56090	=>	6986,
		56091	=>	6988,
		56092	=>	6990,
		56093	=>	6992,
		56094	=>	6993,
		56095	=>	6995,
		56096	=>	6997,
		56097	=>	6999,
		56098	=>	7001,
		56099	=>	7003,
		56100	=>	7005,
		56101	=>	7007,
		56102	=>	7009,
		56103	=>	7011,
		56104	=>	7013,
		56105	=>	7015,
		56106	=>	7017,
		56107	=>	7019,
		56108	=>	7021,
		56109	=>	7023,
		56110	=>	7025,
		56111	=>	7026,
		56112	=>	7028,
		56113	=>	7030,
		56114	=>	7032,
		56115	=>	7034,
		56116	=>	7036,
		56117	=>	7038,
		56118	=>	7040,
		56119	=>	7042,
		56120	=>	7044,
		56121	=>	7046,
		56122	=>	7048,
		56123	=>	7050,
		56124	=>	7052,
		56125	=>	7054,
		56126	=>	7056,
		56127	=>	7058,
		56128	=>	7060,
		56129	=>	7061,
		56130	=>	7063,
		56131	=>	7065,
		56132	=>	7067,
		56133	=>	7069,
		56134	=>	7071,
		56135	=>	7073,
		56136	=>	7075,
		56137	=>	7077,
		56138	=>	7079,
		56139	=>	7081,
		56140	=>	7083,
		56141	=>	7085,
		56142	=>	7087,
		56143	=>	7089,
		56144	=>	7091,
		56145	=>	7093,
		56146	=>	7095,
		56147	=>	7097,
		56148	=>	7099,
		56149	=>	7101,
		56150	=>	7102,
		56151	=>	7104,
		56152	=>	7106,
		56153	=>	7108,
		56154	=>	7110,
		56155	=>	7112,
		56156	=>	7114,
		56157	=>	7116,
		56158	=>	7118,
		56159	=>	7120,
		56160	=>	7122,
		56161	=>	7124,
		56162	=>	7126,
		56163	=>	7128,
		56164	=>	7130,
		56165	=>	7132,
		56166	=>	7134,
		56167	=>	7136,
		56168	=>	7138,
		56169	=>	7140,
		56170	=>	7142,
		56171	=>	7144,
		56172	=>	7145,
		56173	=>	7147,
		56174	=>	7149,
		56175	=>	7151,
		56176	=>	7153,
		56177	=>	7155,
		56178	=>	7157,
		56179	=>	7159,
		56180	=>	7161,
		56181	=>	7163,
		56182	=>	7165,
		56183	=>	7167,
		56184	=>	7169,
		56185	=>	7171,
		56186	=>	7173,
		56187	=>	7175,
		56188	=>	7177,
		56189	=>	7179,
		56190	=>	7181,
		56191	=>	7183,
		56192	=>	7185,
		56193	=>	7187,
		56194	=>	7189,
		56195	=>	7191,
		56196	=>	7193,
		56197	=>	7195,
		56198	=>	7196,
		56199	=>	7198,
		56200	=>	7200,
		56201	=>	7202,
		56202	=>	7204,
		56203	=>	7206,
		56204	=>	7208,
		56205	=>	7210,
		56206	=>	7212,
		56207	=>	7214,
		56208	=>	7216,
		56209	=>	7218,
		56210	=>	7220,
		56211	=>	7222,
		56212	=>	7224,
		56213	=>	7226,
		56214	=>	7228,
		56215	=>	7230,
		56216	=>	7232,
		56217	=>	7234,
		56218	=>	7236,
		56219	=>	7238,
		56220	=>	7240,
		56221	=>	7242,
		56222	=>	7244,
		56223	=>	7246,
		56224	=>	7248,
		56225	=>	7250,
		56226	=>	7252,
		56227	=>	7254,
		56228	=>	7256,
		56229	=>	7257,
		56230	=>	7259,
		56231	=>	7261,
		56232	=>	7263,
		56233	=>	7265,
		56234	=>	7267,
		56235	=>	7269,
		56236	=>	7271,
		56237	=>	7273,
		56238	=>	7275,
		56239	=>	7277,
		56240	=>	7279,
		56241	=>	7281,
		56242	=>	7283,
		56243	=>	7285,
		56244	=>	7287,
		56245	=>	7289,
		56246	=>	7291,
		56247	=>	7293,
		56248	=>	7295,
		56249	=>	7297,
		56250	=>	7299,
		56251	=>	7301,
		56252	=>	7303,
		56253	=>	7305,
		56254	=>	7307,
		56255	=>	7309,
		56256	=>	7311,
		56257	=>	7313,
		56258	=>	7315,
		56259	=>	7317,
		56260	=>	7319,
		56261	=>	7321,
		56262	=>	7323,
		56263	=>	7325,
		56264	=>	7327,
		56265	=>	7329,
		56266	=>	7331,
		56267	=>	7333,
		56268	=>	7335,
		56269	=>	7337,
		56270	=>	7339,
		56271	=>	7341,
		56272	=>	7342,
		56273	=>	7344,
		56274	=>	7346,
		56275	=>	7348,
		56276	=>	7350,
		56277	=>	7352,
		56278	=>	7354,
		56279	=>	7356,
		56280	=>	7358,
		56281	=>	7360,
		56282	=>	7362,
		56283	=>	7364,
		56284	=>	7366,
		56285	=>	7368,
		56286	=>	7370,
		56287	=>	7372,
		56288	=>	7374,
		56289	=>	7376,
		56290	=>	7378,
		56291	=>	7380,
		56292	=>	7382,
		56293	=>	7384,
		56294	=>	7386,
		56295	=>	7388,
		56296	=>	7390,
		56297	=>	7392,
		56298	=>	7394,
		56299	=>	7396,
		56300	=>	7398,
		56301	=>	7400,
		56302	=>	7402,
		56303	=>	7404,
		56304	=>	7406,
		56305	=>	7408,
		56306	=>	7410,
		56307	=>	7412,
		56308	=>	7414,
		56309	=>	7416,
		56310	=>	7418,
		56311	=>	7420,
		56312	=>	7422,
		56313	=>	7424,
		56314	=>	7426,
		56315	=>	7428,
		56316	=>	7430,
		56317	=>	7432,
		56318	=>	7434,
		56319	=>	7436,
		56320	=>	7438,
		56321	=>	7440,
		56322	=>	7442,
		56323	=>	7444,
		56324	=>	7446,
		56325	=>	7448,
		56326	=>	7450,
		56327	=>	7452,
		56328	=>	7454,
		56329	=>	7456,
		56330	=>	7458,
		56331	=>	7460,
		56332	=>	7462,
		56333	=>	7464,
		56334	=>	7466,
		56335	=>	7468,
		56336	=>	7470,
		56337	=>	7472,
		56338	=>	7474,
		56339	=>	7476,
		56340	=>	7478,
		56341	=>	7480,
		56342	=>	7482,
		56343	=>	7484,
		56344	=>	7486,
		56345	=>	7488,
		56346	=>	7490,
		56347	=>	7492,
		56348	=>	7494,
		56349	=>	7496,
		56350	=>	7498,
		56351	=>	7500,
		56352	=>	7502,
		56353	=>	7504,
		56354	=>	7506,
		56355	=>	7508,
		56356	=>	7510,
		56357	=>	7512,
		56358	=>	7514,
		56359	=>	7516,
		56360	=>	7518,
		56361	=>	7520,
		56362	=>	7522,
		56363	=>	7524,
		56364	=>	7526,
		56365	=>	7528,
		56366	=>	7530,
		56367	=>	7532,
		56368	=>	7534,
		56369	=>	7536,
		56370	=>	7538,
		56371	=>	7540,
		56372	=>	7542,
		56373	=>	7544,
		56374	=>	7546,
		56375	=>	7548,
		56376	=>	7550,
		56377	=>	7552,
		56378	=>	7554,
		56379	=>	7556,
		56380	=>	7558,
		56381	=>	7560,
		56382	=>	7562,
		56383	=>	7564,
		56384	=>	7566,
		56385	=>	7568,
		56386	=>	7570,
		56387	=>	7572,
		56388	=>	7574,
		56389	=>	7576,
		56390	=>	7578,
		56391	=>	7580,
		56392	=>	7582,
		56393	=>	7584,
		56394	=>	7586,
		56395	=>	7588,
		56396	=>	7590,
		56397	=>	7592,
		56398	=>	7594,
		56399	=>	7596,
		56400	=>	7598,
		56401	=>	7600,
		56402	=>	7602,
		56403	=>	7604,
		56404	=>	7606,
		56405	=>	7608,
		56406	=>	7610,
		56407	=>	7612,
		56408	=>	7614,
		56409	=>	7616,
		56410	=>	7618,
		56411	=>	7620,
		56412	=>	7622,
		56413	=>	7624,
		56414	=>	7626,
		56415	=>	7628,
		56416	=>	7630,
		56417	=>	7632,
		56418	=>	7634,
		56419	=>	7636,
		56420	=>	7638,
		56421	=>	7640,
		56422	=>	7642,
		56423	=>	7644,
		56424	=>	7646,
		56425	=>	7648,
		56426	=>	7650,
		56427	=>	7652,
		56428	=>	7654,
		56429	=>	7656,
		56430	=>	7659,
		56431	=>	7661,
		56432	=>	7663,
		56433	=>	7665,
		56434	=>	7667,
		56435	=>	7669,
		56436	=>	7671,
		56437	=>	7673,
		56438	=>	7675,
		56439	=>	7677,
		56440	=>	7679,
		56441	=>	7681,
		56442	=>	7683,
		56443	=>	7685,
		56444	=>	7687,
		56445	=>	7689,
		56446	=>	7691,
		56447	=>	7693,
		56448	=>	7695,
		56449	=>	7697,
		56450	=>	7699,
		56451	=>	7701,
		56452	=>	7703,
		56453	=>	7705,
		56454	=>	7707,
		56455	=>	7709,
		56456	=>	7711,
		56457	=>	7713,
		56458	=>	7715,
		56459	=>	7717,
		56460	=>	7719,
		56461	=>	7721,
		56462	=>	7723,
		56463	=>	7725,
		56464	=>	7727,
		56465	=>	7729,
		56466	=>	7731,
		56467	=>	7733,
		56468	=>	7735,
		56469	=>	7737,
		56470	=>	7739,
		56471	=>	7741,
		56472	=>	7743,
		56473	=>	7746,
		56474	=>	7748,
		56475	=>	7750,
		56476	=>	7752,
		56477	=>	7754,
		56478	=>	7756,
		56479	=>	7758,
		56480	=>	7760,
		56481	=>	7762,
		56482	=>	7764,
		56483	=>	7766,
		56484	=>	7768,
		56485	=>	7770,
		56486	=>	7772,
		56487	=>	7774,
		56488	=>	7776,
		56489	=>	7778,
		56490	=>	7780,
		56491	=>	7782,
		56492	=>	7784,
		56493	=>	7786,
		56494	=>	7788,
		56495	=>	7790,
		56496	=>	7792,
		56497	=>	7794,
		56498	=>	7796,
		56499	=>	7798,
		56500	=>	7800,
		56501	=>	7802,
		56502	=>	7804,
		56503	=>	7806,
		56504	=>	7809,
		56505	=>	7811,
		56506	=>	7813,
		56507	=>	7815,
		56508	=>	7817,
		56509	=>	7819,
		56510	=>	7821,
		56511	=>	7823,
		56512	=>	7825,
		56513	=>	7827,
		56514	=>	7829,
		56515	=>	7831,
		56516	=>	7833,
		56517	=>	7835,
		56518	=>	7837,
		56519	=>	7839,
		56520	=>	7841,
		56521	=>	7843,
		56522	=>	7845,
		56523	=>	7847,
		56524	=>	7849,
		56525	=>	7851,
		56526	=>	7853,
		56527	=>	7855,
		56528	=>	7857,
		56529	=>	7859,
		56530	=>	7862,
		56531	=>	7864,
		56532	=>	7866,
		56533	=>	7868,
		56534	=>	7870,
		56535	=>	7872,
		56536	=>	7874,
		56537	=>	7876,
		56538	=>	7878,
		56539	=>	7880,
		56540	=>	7882,
		56541	=>	7884,
		56542	=>	7886,
		56543	=>	7888,
		56544	=>	7890,
		56545	=>	7892,
		56546	=>	7894,
		56547	=>	7896,
		56548	=>	7898,
		56549	=>	7900,
		56550	=>	7902,
		56551	=>	7904,
		56552	=>	7906,
		56553	=>	7909,
		56554	=>	7911,
		56555	=>	7913,
		56556	=>	7915,
		56557	=>	7917,
		56558	=>	7919,
		56559	=>	7921,
		56560	=>	7923,
		56561	=>	7925,
		56562	=>	7927,
		56563	=>	7929,
		56564	=>	7931,
		56565	=>	7933,
		56566	=>	7935,
		56567	=>	7937,
		56568	=>	7939,
		56569	=>	7941,
		56570	=>	7943,
		56571	=>	7945,
		56572	=>	7947,
		56573	=>	7950,
		56574	=>	7952,
		56575	=>	7954,
		56576	=>	7956,
		56577	=>	7958,
		56578	=>	7960,
		56579	=>	7962,
		56580	=>	7964,
		56581	=>	7966,
		56582	=>	7968,
		56583	=>	7970,
		56584	=>	7972,
		56585	=>	7974,
		56586	=>	7976,
		56587	=>	7978,
		56588	=>	7980,
		56589	=>	7982,
		56590	=>	7984,
		56591	=>	7986,
		56592	=>	7989,
		56593	=>	7991,
		56594	=>	7993,
		56595	=>	7995,
		56596	=>	7997,
		56597	=>	7999,
		56598	=>	8001,
		56599	=>	8003,
		56600	=>	8005,
		56601	=>	8007,
		56602	=>	8009,
		56603	=>	8011,
		56604	=>	8013,
		56605	=>	8015,
		56606	=>	8017,
		56607	=>	8019,
		56608	=>	8021,
		56609	=>	8023,
		56610	=>	8026,
		56611	=>	8028,
		56612	=>	8030,
		56613	=>	8032,
		56614	=>	8034,
		56615	=>	8036,
		56616	=>	8038,
		56617	=>	8040,
		56618	=>	8042,
		56619	=>	8044,
		56620	=>	8046,
		56621	=>	8048,
		56622	=>	8050,
		56623	=>	8052,
		56624	=>	8054,
		56625	=>	8056,
		56626	=>	8059,
		56627	=>	8061,
		56628	=>	8063,
		56629	=>	8065,
		56630	=>	8067,
		56631	=>	8069,
		56632	=>	8071,
		56633	=>	8073,
		56634	=>	8075,
		56635	=>	8077,
		56636	=>	8079,
		56637	=>	8081,
		56638	=>	8083,
		56639	=>	8085,
		56640	=>	8087,
		56641	=>	8090,
		56642	=>	8092,
		56643	=>	8094,
		56644	=>	8096,
		56645	=>	8098,
		56646	=>	8100,
		56647	=>	8102,
		56648	=>	8104,
		56649	=>	8106,
		56650	=>	8108,
		56651	=>	8110,
		56652	=>	8112,
		56653	=>	8114,
		56654	=>	8116,
		56655	=>	8118,
		56656	=>	8121,
		56657	=>	8123,
		56658	=>	8125,
		56659	=>	8127,
		56660	=>	8129,
		56661	=>	8131,
		56662	=>	8133,
		56663	=>	8135,
		56664	=>	8137,
		56665	=>	8139,
		56666	=>	8141,
		56667	=>	8143,
		56668	=>	8145,
		56669	=>	8147,
		56670	=>	8150,
		56671	=>	8152,
		56672	=>	8154,
		56673	=>	8156,
		56674	=>	8158,
		56675	=>	8160,
		56676	=>	8162,
		56677	=>	8164,
		56678	=>	8166,
		56679	=>	8168,
		56680	=>	8170,
		56681	=>	8172,
		56682	=>	8174,
		56683	=>	8177,
		56684	=>	8179,
		56685	=>	8181,
		56686	=>	8183,
		56687	=>	8185,
		56688	=>	8187,
		56689	=>	8189,
		56690	=>	8191,
		56691	=>	8193,
		56692	=>	8195,
		56693	=>	8197,
		56694	=>	8199,
		56695	=>	8201,
		56696	=>	8204,
		56697	=>	8206,
		56698	=>	8208,
		56699	=>	8210,
		56700	=>	8212,
		56701	=>	8214,
		56702	=>	8216,
		56703	=>	8218,
		56704	=>	8220,
		56705	=>	8222,
		56706	=>	8224,
		56707	=>	8226,
		56708	=>	8228,
		56709	=>	8231,
		56710	=>	8233,
		56711	=>	8235,
		56712	=>	8237,
		56713	=>	8239,
		56714	=>	8241,
		56715	=>	8243,
		56716	=>	8245,
		56717	=>	8247,
		56718	=>	8249,
		56719	=>	8251,
		56720	=>	8253,
		56721	=>	8256,
		56722	=>	8258,
		56723	=>	8260,
		56724	=>	8262,
		56725	=>	8264,
		56726	=>	8266,
		56727	=>	8268,
		56728	=>	8270,
		56729	=>	8272,
		56730	=>	8274,
		56731	=>	8276,
		56732	=>	8279,
		56733	=>	8281,
		56734	=>	8283,
		56735	=>	8285,
		56736	=>	8287,
		56737	=>	8289,
		56738	=>	8291,
		56739	=>	8293,
		56740	=>	8295,
		56741	=>	8297,
		56742	=>	8299,
		56743	=>	8302,
		56744	=>	8304,
		56745	=>	8306,
		56746	=>	8308,
		56747	=>	8310,
		56748	=>	8312,
		56749	=>	8314,
		56750	=>	8316,
		56751	=>	8318,
		56752	=>	8320,
		56753	=>	8322,
		56754	=>	8325,
		56755	=>	8327,
		56756	=>	8329,
		56757	=>	8331,
		56758	=>	8333,
		56759	=>	8335,
		56760	=>	8337,
		56761	=>	8339,
		56762	=>	8341,
		56763	=>	8343,
		56764	=>	8345,
		56765	=>	8348,
		56766	=>	8350,
		56767	=>	8352,
		56768	=>	8354,
		56769	=>	8356,
		56770	=>	8358,
		56771	=>	8360,
		56772	=>	8362,
		56773	=>	8364,
		56774	=>	8366,
		56775	=>	8368,
		56776	=>	8371,
		56777	=>	8373,
		56778	=>	8375,
		56779	=>	8377,
		56780	=>	8379,
		56781	=>	8381,
		56782	=>	8383,
		56783	=>	8385,
		56784	=>	8387,
		56785	=>	8389,
		56786	=>	8392,
		56787	=>	8394,
		56788	=>	8396,
		56789	=>	8398,
		56790	=>	8400,
		56791	=>	8402,
		56792	=>	8404,
		56793	=>	8406,
		56794	=>	8408,
		56795	=>	8410,
		56796	=>	8413,
		56797	=>	8415,
		56798	=>	8417,
		56799	=>	8419,
		56800	=>	8421,
		56801	=>	8423,
		56802	=>	8425,
		56803	=>	8427,
		56804	=>	8429,
		56805	=>	8432,
		56806	=>	8434,
		56807	=>	8436,
		56808	=>	8438,
		56809	=>	8440,
		56810	=>	8442,
		56811	=>	8444,
		56812	=>	8446,
		56813	=>	8448,
		56814	=>	8450,
		56815	=>	8453,
		56816	=>	8455,
		56817	=>	8457,
		56818	=>	8459,
		56819	=>	8461,
		56820	=>	8463,
		56821	=>	8465,
		56822	=>	8467,
		56823	=>	8469,
		56824	=>	8472,
		56825	=>	8474,
		56826	=>	8476,
		56827	=>	8478,
		56828	=>	8480,
		56829	=>	8482,
		56830	=>	8484,
		56831	=>	8486,
		56832	=>	8488,
		56833	=>	8490,
		56834	=>	8493,
		56835	=>	8495,
		56836	=>	8497,
		56837	=>	8499,
		56838	=>	8501,
		56839	=>	8503,
		56840	=>	8505,
		56841	=>	8507,
		56842	=>	8509,
		56843	=>	8512,
		56844	=>	8514,
		56845	=>	8516,
		56846	=>	8518,
		56847	=>	8520,
		56848	=>	8522,
		56849	=>	8524,
		56850	=>	8526,
		56851	=>	8529,
		56852	=>	8531,
		56853	=>	8533,
		56854	=>	8535,
		56855	=>	8537,
		56856	=>	8539,
		56857	=>	8541,
		56858	=>	8543,
		56859	=>	8545,
		56860	=>	8548,
		56861	=>	8550,
		56862	=>	8552,
		56863	=>	8554,
		56864	=>	8556,
		56865	=>	8558,
		56866	=>	8560,
		56867	=>	8562,
		56868	=>	8564,
		56869	=>	8567,
		56870	=>	8569,
		56871	=>	8571,
		56872	=>	8573,
		56873	=>	8575,
		56874	=>	8577,
		56875	=>	8579,
		56876	=>	8581,
		56877	=>	8584,
		56878	=>	8586,
		56879	=>	8588,
		56880	=>	8590,
		56881	=>	8592,
		56882	=>	8594,
		56883	=>	8596,
		56884	=>	8598,
		56885	=>	8601,
		56886	=>	8603,
		56887	=>	8605,
		56888	=>	8607,
		56889	=>	8609,
		56890	=>	8611,
		56891	=>	8613,
		56892	=>	8615,
		56893	=>	8617,
		56894	=>	8620,
		56895	=>	8622,
		56896	=>	8624,
		56897	=>	8626,
		56898	=>	8628,
		56899	=>	8630,
		56900	=>	8632,
		56901	=>	8634,
		56902	=>	8637,
		56903	=>	8639,
		56904	=>	8641,
		56905	=>	8643,
		56906	=>	8645,
		56907	=>	8647,
		56908	=>	8649,
		56909	=>	8651,
		56910	=>	8654,
		56911	=>	8656,
		56912	=>	8658,
		56913	=>	8660,
		56914	=>	8662,
		56915	=>	8664,
		56916	=>	8666,
		56917	=>	8669,
		56918	=>	8671,
		56919	=>	8673,
		56920	=>	8675,
		56921	=>	8677,
		56922	=>	8679,
		56923	=>	8681,
		56924	=>	8683,
		56925	=>	8686,
		56926	=>	8688,
		56927	=>	8690,
		56928	=>	8692,
		56929	=>	8694,
		56930	=>	8696,
		56931	=>	8698,
		56932	=>	8700,
		56933	=>	8703,
		56934	=>	8705,
		56935	=>	8707,
		56936	=>	8709,
		56937	=>	8711,
		56938	=>	8713,
		56939	=>	8715,
		56940	=>	8718,
		56941	=>	8720,
		56942	=>	8722,
		56943	=>	8724,
		56944	=>	8726,
		56945	=>	8728,
		56946	=>	8730,
		56947	=>	8732,
		56948	=>	8735,
		56949	=>	8737,
		56950	=>	8739,
		56951	=>	8741,
		56952	=>	8743,
		56953	=>	8745,
		56954	=>	8747,
		56955	=>	8750,
		56956	=>	8752,
		56957	=>	8754,
		56958	=>	8756,
		56959	=>	8758,
		56960	=>	8760,
		56961	=>	8762,
		56962	=>	8765,
		56963	=>	8767,
		56964	=>	8769,
		56965	=>	8771,
		56966	=>	8773,
		56967	=>	8775,
		56968	=>	8777,
		56969	=>	8780,
		56970	=>	8782,
		56971	=>	8784,
		56972	=>	8786,
		56973	=>	8788,
		56974	=>	8790,
		56975	=>	8792,
		56976	=>	8794,
		56977	=>	8797,
		56978	=>	8799,
		56979	=>	8801,
		56980	=>	8803,
		56981	=>	8805,
		56982	=>	8807,
		56983	=>	8809,
		56984	=>	8812,
		56985	=>	8814,
		56986	=>	8816,
		56987	=>	8818,
		56988	=>	8820,
		56989	=>	8822,
		56990	=>	8824,
		56991	=>	8827,
		56992	=>	8829,
		56993	=>	8831,
		56994	=>	8833,
		56995	=>	8835,
		56996	=>	8837,
		56997	=>	8840,
		56998	=>	8842,
		56999	=>	8844,
		57000	=>	8846,
		57001	=>	8848,
		57002	=>	8850,
		57003	=>	8852,
		57004	=>	8855,
		57005	=>	8857,
		57006	=>	8859,
		57007	=>	8861,
		57008	=>	8863,
		57009	=>	8865,
		57010	=>	8867,
		57011	=>	8870,
		57012	=>	8872,
		57013	=>	8874,
		57014	=>	8876,
		57015	=>	8878,
		57016	=>	8880,
		57017	=>	8882,
		57018	=>	8885,
		57019	=>	8887,
		57020	=>	8889,
		57021	=>	8891,
		57022	=>	8893,
		57023	=>	8895,
		57024	=>	8898,
		57025	=>	8900,
		57026	=>	8902,
		57027	=>	8904,
		57028	=>	8906,
		57029	=>	8908,
		57030	=>	8910,
		57031	=>	8913,
		57032	=>	8915,
		57033	=>	8917,
		57034	=>	8919,
		57035	=>	8921,
		57036	=>	8923,
		57037	=>	8926,
		57038	=>	8928,
		57039	=>	8930,
		57040	=>	8932,
		57041	=>	8934,
		57042	=>	8936,
		57043	=>	8938,
		57044	=>	8941,
		57045	=>	8943,
		57046	=>	8945,
		57047	=>	8947,
		57048	=>	8949,
		57049	=>	8951,
		57050	=>	8954,
		57051	=>	8956,
		57052	=>	8958,
		57053	=>	8960,
		57054	=>	8962,
		57055	=>	8964,
		57056	=>	8967,
		57057	=>	8969,
		57058	=>	8971,
		57059	=>	8973,
		57060	=>	8975,
		57061	=>	8977,
		57062	=>	8979,
		57063	=>	8982,
		57064	=>	8984,
		57065	=>	8986,
		57066	=>	8988,
		57067	=>	8990,
		57068	=>	8992,
		57069	=>	8995,
		57070	=>	8997,
		57071	=>	8999,
		57072	=>	9001,
		57073	=>	9003,
		57074	=>	9005,
		57075	=>	9008,
		57076	=>	9010,
		57077	=>	9012,
		57078	=>	9014,
		57079	=>	9016,
		57080	=>	9018,
		57081	=>	9021,
		57082	=>	9023,
		57083	=>	9025,
		57084	=>	9027,
		57085	=>	9029,
		57086	=>	9031,
		57087	=>	9034,
		57088	=>	9036,
		57089	=>	9038,
		57090	=>	9040,
		57091	=>	9042,
		57092	=>	9044,
		57093	=>	9047,
		57094	=>	9049,
		57095	=>	9051,
		57096	=>	9053,
		57097	=>	9055,
		57098	=>	9057,
		57099	=>	9060,
		57100	=>	9062,
		57101	=>	9064,
		57102	=>	9066,
		57103	=>	9068,
		57104	=>	9070,
		57105	=>	9073,
		57106	=>	9075,
		57107	=>	9077,
		57108	=>	9079,
		57109	=>	9081,
		57110	=>	9083,
		57111	=>	9086,
		57112	=>	9088,
		57113	=>	9090,
		57114	=>	9092,
		57115	=>	9094,
		57116	=>	9096,
		57117	=>	9099,
		57118	=>	9101,
		57119	=>	9103,
		57120	=>	9105,
		57121	=>	9107,
		57122	=>	9110,
		57123	=>	9112,
		57124	=>	9114,
		57125	=>	9116,
		57126	=>	9118,
		57127	=>	9120,
		57128	=>	9123,
		57129	=>	9125,
		57130	=>	9127,
		57131	=>	9129,
		57132	=>	9131,
		57133	=>	9133,
		57134	=>	9136,
		57135	=>	9138,
		57136	=>	9140,
		57137	=>	9142,
		57138	=>	9144,
		57139	=>	9146,
		57140	=>	9149,
		57141	=>	9151,
		57142	=>	9153,
		57143	=>	9155,
		57144	=>	9157,
		57145	=>	9160,
		57146	=>	9162,
		57147	=>	9164,
		57148	=>	9166,
		57149	=>	9168,
		57150	=>	9170,
		57151	=>	9173,
		57152	=>	9175,
		57153	=>	9177,
		57154	=>	9179,
		57155	=>	9181,
		57156	=>	9184,
		57157	=>	9186,
		57158	=>	9188,
		57159	=>	9190,
		57160	=>	9192,
		57161	=>	9194,
		57162	=>	9197,
		57163	=>	9199,
		57164	=>	9201,
		57165	=>	9203,
		57166	=>	9205,
		57167	=>	9208,
		57168	=>	9210,
		57169	=>	9212,
		57170	=>	9214,
		57171	=>	9216,
		57172	=>	9218,
		57173	=>	9221,
		57174	=>	9223,
		57175	=>	9225,
		57176	=>	9227,
		57177	=>	9229,
		57178	=>	9232,
		57179	=>	9234,
		57180	=>	9236,
		57181	=>	9238,
		57182	=>	9240,
		57183	=>	9243,
		57184	=>	9245,
		57185	=>	9247,
		57186	=>	9249,
		57187	=>	9251,
		57188	=>	9253,
		57189	=>	9256,
		57190	=>	9258,
		57191	=>	9260,
		57192	=>	9262,
		57193	=>	9264,
		57194	=>	9267,
		57195	=>	9269,
		57196	=>	9271,
		57197	=>	9273,
		57198	=>	9275,
		57199	=>	9278,
		57200	=>	9280,
		57201	=>	9282,
		57202	=>	9284,
		57203	=>	9286,
		57204	=>	9288,
		57205	=>	9291,
		57206	=>	9293,
		57207	=>	9295,
		57208	=>	9297,
		57209	=>	9299,
		57210	=>	9302,
		57211	=>	9304,
		57212	=>	9306,
		57213	=>	9308,
		57214	=>	9310,
		57215	=>	9313,
		57216	=>	9315,
		57217	=>	9317,
		57218	=>	9319,
		57219	=>	9321,
		57220	=>	9324,
		57221	=>	9326,
		57222	=>	9328,
		57223	=>	9330,
		57224	=>	9332,
		57225	=>	9335,
		57226	=>	9337,
		57227	=>	9339,
		57228	=>	9341,
		57229	=>	9343,
		57230	=>	9346,
		57231	=>	9348,
		57232	=>	9350,
		57233	=>	9352,
		57234	=>	9354,
		57235	=>	9357,
		57236	=>	9359,
		57237	=>	9361,
		57238	=>	9363,
		57239	=>	9365,
		57240	=>	9368,
		57241	=>	9370,
		57242	=>	9372,
		57243	=>	9374,
		57244	=>	9376,
		57245	=>	9379,
		57246	=>	9381,
		57247	=>	9383,
		57248	=>	9385,
		57249	=>	9387,
		57250	=>	9390,
		57251	=>	9392,
		57252	=>	9394,
		57253	=>	9396,
		57254	=>	9398,
		57255	=>	9401,
		57256	=>	9403,
		57257	=>	9405,
		57258	=>	9407,
		57259	=>	9409,
		57260	=>	9412,
		57261	=>	9414,
		57262	=>	9416,
		57263	=>	9418,
		57264	=>	9420,
		57265	=>	9423,
		57266	=>	9425,
		57267	=>	9427,
		57268	=>	9429,
		57269	=>	9431,
		57270	=>	9434,
		57271	=>	9436,
		57272	=>	9438,
		57273	=>	9440,
		57274	=>	9442,
		57275	=>	9445,
		57276	=>	9447,
		57277	=>	9449,
		57278	=>	9451,
		57279	=>	9453,
		57280	=>	9456,
		57281	=>	9458,
		57282	=>	9460,
		57283	=>	9462,
		57284	=>	9464,
		57285	=>	9467,
		57286	=>	9469,
		57287	=>	9471,
		57288	=>	9473,
		57289	=>	9476,
		57290	=>	9478,
		57291	=>	9480,
		57292	=>	9482,
		57293	=>	9484,
		57294	=>	9487,
		57295	=>	9489,
		57296	=>	9491,
		57297	=>	9493,
		57298	=>	9495,
		57299	=>	9498,
		57300	=>	9500,
		57301	=>	9502,
		57302	=>	9504,
		57303	=>	9506,
		57304	=>	9509,
		57305	=>	9511,
		57306	=>	9513,
		57307	=>	9515,
		57308	=>	9518,
		57309	=>	9520,
		57310	=>	9522,
		57311	=>	9524,
		57312	=>	9526,
		57313	=>	9529,
		57314	=>	9531,
		57315	=>	9533,
		57316	=>	9535,
		57317	=>	9537,
		57318	=>	9540,
		57319	=>	9542,
		57320	=>	9544,
		57321	=>	9546,
		57322	=>	9549,
		57323	=>	9551,
		57324	=>	9553,
		57325	=>	9555,
		57326	=>	9557,
		57327	=>	9560,
		57328	=>	9562,
		57329	=>	9564,
		57330	=>	9566,
		57331	=>	9569,
		57332	=>	9571,
		57333	=>	9573,
		57334	=>	9575,
		57335	=>	9577,
		57336	=>	9580,
		57337	=>	9582,
		57338	=>	9584,
		57339	=>	9586,
		57340	=>	9588,
		57341	=>	9591,
		57342	=>	9593,
		57343	=>	9595,
		57344	=>	9597,
		57345	=>	9600,
		57346	=>	9602,
		57347	=>	9604,
		57348	=>	9606,
		57349	=>	9608,
		57350	=>	9611,
		57351	=>	9613,
		57352	=>	9615,
		57353	=>	9617,
		57354	=>	9620,
		57355	=>	9622,
		57356	=>	9624,
		57357	=>	9626,
		57358	=>	9628,
		57359	=>	9631,
		57360	=>	9633,
		57361	=>	9635,
		57362	=>	9637,
		57363	=>	9640,
		57364	=>	9642,
		57365	=>	9644,
		57366	=>	9646,
		57367	=>	9649,
		57368	=>	9651,
		57369	=>	9653,
		57370	=>	9655,
		57371	=>	9657,
		57372	=>	9660,
		57373	=>	9662,
		57374	=>	9664,
		57375	=>	9666,
		57376	=>	9669,
		57377	=>	9671,
		57378	=>	9673,
		57379	=>	9675,
		57380	=>	9677,
		57381	=>	9680,
		57382	=>	9682,
		57383	=>	9684,
		57384	=>	9686,
		57385	=>	9689,
		57386	=>	9691,
		57387	=>	9693,
		57388	=>	9695,
		57389	=>	9698,
		57390	=>	9700,
		57391	=>	9702,
		57392	=>	9704,
		57393	=>	9706,
		57394	=>	9709,
		57395	=>	9711,
		57396	=>	9713,
		57397	=>	9715,
		57398	=>	9718,
		57399	=>	9720,
		57400	=>	9722,
		57401	=>	9724,
		57402	=>	9727,
		57403	=>	9729,
		57404	=>	9731,
		57405	=>	9733,
		57406	=>	9736,
		57407	=>	9738,
		57408	=>	9740,
		57409	=>	9742,
		57410	=>	9744,
		57411	=>	9747,
		57412	=>	9749,
		57413	=>	9751,
		57414	=>	9753,
		57415	=>	9756,
		57416	=>	9758,
		57417	=>	9760,
		57418	=>	9762,
		57419	=>	9765,
		57420	=>	9767,
		57421	=>	9769,
		57422	=>	9771,
		57423	=>	9774,
		57424	=>	9776,
		57425	=>	9778,
		57426	=>	9780,
		57427	=>	9782,
		57428	=>	9785,
		57429	=>	9787,
		57430	=>	9789,
		57431	=>	9791,
		57432	=>	9794,
		57433	=>	9796,
		57434	=>	9798,
		57435	=>	9800,
		57436	=>	9803,
		57437	=>	9805,
		57438	=>	9807,
		57439	=>	9809,
		57440	=>	9812,
		57441	=>	9814,
		57442	=>	9816,
		57443	=>	9818,
		57444	=>	9821,
		57445	=>	9823,
		57446	=>	9825,
		57447	=>	9827,
		57448	=>	9830,
		57449	=>	9832,
		57450	=>	9834,
		57451	=>	9836,
		57452	=>	9839,
		57453	=>	9841,
		57454	=>	9843,
		57455	=>	9845,
		57456	=>	9848,
		57457	=>	9850,
		57458	=>	9852,
		57459	=>	9854,
		57460	=>	9856,
		57461	=>	9859,
		57462	=>	9861,
		57463	=>	9863,
		57464	=>	9865,
		57465	=>	9868,
		57466	=>	9870,
		57467	=>	9872,
		57468	=>	9874,
		57469	=>	9877,
		57470	=>	9879,
		57471	=>	9881,
		57472	=>	9883,
		57473	=>	9886,
		57474	=>	9888,
		57475	=>	9890,
		57476	=>	9892,
		57477	=>	9895,
		57478	=>	9897,
		57479	=>	9899,
		57480	=>	9901,
		57481	=>	9904,
		57482	=>	9906,
		57483	=>	9908,
		57484	=>	9910,
		57485	=>	9913,
		57486	=>	9915,
		57487	=>	9917,
		57488	=>	9919,
		57489	=>	9922,
		57490	=>	9924,
		57491	=>	9926,
		57492	=>	9928,
		57493	=>	9931,
		57494	=>	9933,
		57495	=>	9935,
		57496	=>	9937,
		57497	=>	9940,
		57498	=>	9942,
		57499	=>	9944,
		57500	=>	9946,
		57501	=>	9949,
		57502	=>	9951,
		57503	=>	9953,
		57504	=>	9956,
		57505	=>	9958,
		57506	=>	9960,
		57507	=>	9962,
		57508	=>	9965,
		57509	=>	9967,
		57510	=>	9969,
		57511	=>	9971,
		57512	=>	9974,
		57513	=>	9976,
		57514	=>	9978,
		57515	=>	9980,
		57516	=>	9983,
		57517	=>	9985,
		57518	=>	9987,
		57519	=>	9989,
		57520	=>	9992,
		57521	=>	9994,
		57522	=>	9996,
		57523	=>	9998,
		57524	=>	10001,
		57525	=>	10003,
		57526	=>	10005,
		57527	=>	10007,
		57528	=>	10010,
		57529	=>	10012,
		57530	=>	10014,
		57531	=>	10016,
		57532	=>	10019,
		57533	=>	10021,
		57534	=>	10023,
		57535	=>	10026,
		57536	=>	10028,
		57537	=>	10030,
		57538	=>	10032,
		57539	=>	10035,
		57540	=>	10037,
		57541	=>	10039,
		57542	=>	10041,
		57543	=>	10044,
		57544	=>	10046,
		57545	=>	10048,
		57546	=>	10050,
		57547	=>	10053,
		57548	=>	10055,
		57549	=>	10057,
		57550	=>	10059,
		57551	=>	10062,
		57552	=>	10064,
		57553	=>	10066,
		57554	=>	10069,
		57555	=>	10071,
		57556	=>	10073,
		57557	=>	10075,
		57558	=>	10078,
		57559	=>	10080,
		57560	=>	10082,
		57561	=>	10084,
		57562	=>	10087,
		57563	=>	10089,
		57564	=>	10091,
		57565	=>	10093,
		57566	=>	10096,
		57567	=>	10098,
		57568	=>	10100,
		57569	=>	10103,
		57570	=>	10105,
		57571	=>	10107,
		57572	=>	10109,
		57573	=>	10112,
		57574	=>	10114,
		57575	=>	10116,
		57576	=>	10118,
		57577	=>	10121,
		57578	=>	10123,
		57579	=>	10125,
		57580	=>	10128,
		57581	=>	10130,
		57582	=>	10132,
		57583	=>	10134,
		57584	=>	10137,
		57585	=>	10139,
		57586	=>	10141,
		57587	=>	10143,
		57588	=>	10146,
		57589	=>	10148,
		57590	=>	10150,
		57591	=>	10153,
		57592	=>	10155,
		57593	=>	10157,
		57594	=>	10159,
		57595	=>	10162,
		57596	=>	10164,
		57597	=>	10166,
		57598	=>	10168,
		57599	=>	10171,
		57600	=>	10173,
		57601	=>	10175,
		57602	=>	10178,
		57603	=>	10180,
		57604	=>	10182,
		57605	=>	10184,
		57606	=>	10187,
		57607	=>	10189,
		57608	=>	10191,
		57609	=>	10193,
		57610	=>	10196,
		57611	=>	10198,
		57612	=>	10200,
		57613	=>	10203,
		57614	=>	10205,
		57615	=>	10207,
		57616	=>	10209,
		57617	=>	10212,
		57618	=>	10214,
		57619	=>	10216,
		57620	=>	10219,
		57621	=>	10221,
		57622	=>	10223,
		57623	=>	10225,
		57624	=>	10228,
		57625	=>	10230,
		57626	=>	10232,
		57627	=>	10234,
		57628	=>	10237,
		57629	=>	10239,
		57630	=>	10241,
		57631	=>	10244,
		57632	=>	10246,
		57633	=>	10248,
		57634	=>	10250,
		57635	=>	10253,
		57636	=>	10255,
		57637	=>	10257,
		57638	=>	10260,
		57639	=>	10262,
		57640	=>	10264,
		57641	=>	10266,
		57642	=>	10269,
		57643	=>	10271,
		57644	=>	10273,
		57645	=>	10276,
		57646	=>	10278,
		57647	=>	10280,
		57648	=>	10282,
		57649	=>	10285,
		57650	=>	10287,
		57651	=>	10289,
		57652	=>	10292,
		57653	=>	10294,
		57654	=>	10296,
		57655	=>	10298,
		57656	=>	10301,
		57657	=>	10303,
		57658	=>	10305,
		57659	=>	10308,
		57660	=>	10310,
		57661	=>	10312,
		57662	=>	10314,
		57663	=>	10317,
		57664	=>	10319,
		57665	=>	10321,
		57666	=>	10324,
		57667	=>	10326,
		57668	=>	10328,
		57669	=>	10330,
		57670	=>	10333,
		57671	=>	10335,
		57672	=>	10337,
		57673	=>	10340,
		57674	=>	10342,
		57675	=>	10344,
		57676	=>	10346,
		57677	=>	10349,
		57678	=>	10351,
		57679	=>	10353,
		57680	=>	10356,
		57681	=>	10358,
		57682	=>	10360,
		57683	=>	10363,
		57684	=>	10365,
		57685	=>	10367,
		57686	=>	10369,
		57687	=>	10372,
		57688	=>	10374,
		57689	=>	10376,
		57690	=>	10379,
		57691	=>	10381,
		57692	=>	10383,
		57693	=>	10385,
		57694	=>	10388,
		57695	=>	10390,
		57696	=>	10392,
		57697	=>	10395,
		57698	=>	10397,
		57699	=>	10399,
		57700	=>	10402,
		57701	=>	10404,
		57702	=>	10406,
		57703	=>	10408,
		57704	=>	10411,
		57705	=>	10413,
		57706	=>	10415,
		57707	=>	10418,
		57708	=>	10420,
		57709	=>	10422,
		57710	=>	10425,
		57711	=>	10427,
		57712	=>	10429,
		57713	=>	10431,
		57714	=>	10434,
		57715	=>	10436,
		57716	=>	10438,
		57717	=>	10441,
		57718	=>	10443,
		57719	=>	10445,
		57720	=>	10448,
		57721	=>	10450,
		57722	=>	10452,
		57723	=>	10454,
		57724	=>	10457,
		57725	=>	10459,
		57726	=>	10461,
		57727	=>	10464,
		57728	=>	10466,
		57729	=>	10468,
		57730	=>	10471,
		57731	=>	10473,
		57732	=>	10475,
		57733	=>	10477,
		57734	=>	10480,
		57735	=>	10482,
		57736	=>	10484,
		57737	=>	10487,
		57738	=>	10489,
		57739	=>	10491,
		57740	=>	10494,
		57741	=>	10496,
		57742	=>	10498,
		57743	=>	10500,
		57744	=>	10503,
		57745	=>	10505,
		57746	=>	10507,
		57747	=>	10510,
		57748	=>	10512,
		57749	=>	10514,
		57750	=>	10517,
		57751	=>	10519,
		57752	=>	10521,
		57753	=>	10524,
		57754	=>	10526,
		57755	=>	10528,
		57756	=>	10530,
		57757	=>	10533,
		57758	=>	10535,
		57759	=>	10537,
		57760	=>	10540,
		57761	=>	10542,
		57762	=>	10544,
		57763	=>	10547,
		57764	=>	10549,
		57765	=>	10551,
		57766	=>	10554,
		57767	=>	10556,
		57768	=>	10558,
		57769	=>	10560,
		57770	=>	10563,
		57771	=>	10565,
		57772	=>	10567,
		57773	=>	10570,
		57774	=>	10572,
		57775	=>	10574,
		57776	=>	10577,
		57777	=>	10579,
		57778	=>	10581,
		57779	=>	10584,
		57780	=>	10586,
		57781	=>	10588,
		57782	=>	10590,
		57783	=>	10593,
		57784	=>	10595,
		57785	=>	10597,
		57786	=>	10600,
		57787	=>	10602,
		57788	=>	10604,
		57789	=>	10607,
		57790	=>	10609,
		57791	=>	10611,
		57792	=>	10614,
		57793	=>	10616,
		57794	=>	10618,
		57795	=>	10621,
		57796	=>	10623,
		57797	=>	10625,
		57798	=>	10628,
		57799	=>	10630,
		57800	=>	10632,
		57801	=>	10634,
		57802	=>	10637,
		57803	=>	10639,
		57804	=>	10641,
		57805	=>	10644,
		57806	=>	10646,
		57807	=>	10648,
		57808	=>	10651,
		57809	=>	10653,
		57810	=>	10655,
		57811	=>	10658,
		57812	=>	10660,
		57813	=>	10662,
		57814	=>	10665,
		57815	=>	10667,
		57816	=>	10669,
		57817	=>	10672,
		57818	=>	10674,
		57819	=>	10676,
		57820	=>	10679,
		57821	=>	10681,
		57822	=>	10683,
		57823	=>	10685,
		57824	=>	10688,
		57825	=>	10690,
		57826	=>	10692,
		57827	=>	10695,
		57828	=>	10697,
		57829	=>	10699,
		57830	=>	10702,
		57831	=>	10704,
		57832	=>	10706,
		57833	=>	10709,
		57834	=>	10711,
		57835	=>	10713,
		57836	=>	10716,
		57837	=>	10718,
		57838	=>	10720,
		57839	=>	10723,
		57840	=>	10725,
		57841	=>	10727,
		57842	=>	10730,
		57843	=>	10732,
		57844	=>	10734,
		57845	=>	10737,
		57846	=>	10739,
		57847	=>	10741,
		57848	=>	10744,
		57849	=>	10746,
		57850	=>	10748,
		57851	=>	10751,
		57852	=>	10753,
		57853	=>	10755,
		57854	=>	10758,
		57855	=>	10760,
		57856	=>	10762,
		57857	=>	10765,
		57858	=>	10767,
		57859	=>	10769,
		57860	=>	10772,
		57861	=>	10774,
		57862	=>	10776,
		57863	=>	10778,
		57864	=>	10781,
		57865	=>	10783,
		57866	=>	10785,
		57867	=>	10788,
		57868	=>	10790,
		57869	=>	10792,
		57870	=>	10795,
		57871	=>	10797,
		57872	=>	10799,
		57873	=>	10802,
		57874	=>	10804,
		57875	=>	10806,
		57876	=>	10809,
		57877	=>	10811,
		57878	=>	10813,
		57879	=>	10816,
		57880	=>	10818,
		57881	=>	10820,
		57882	=>	10823,
		57883	=>	10825,
		57884	=>	10827,
		57885	=>	10830,
		57886	=>	10832,
		57887	=>	10834,
		57888	=>	10837,
		57889	=>	10839,
		57890	=>	10841,
		57891	=>	10844,
		57892	=>	10846,
		57893	=>	10848,
		57894	=>	10851,
		57895	=>	10853,
		57896	=>	10855,
		57897	=>	10858,
		57898	=>	10860,
		57899	=>	10862,
		57900	=>	10865,
		57901	=>	10867,
		57902	=>	10869,
		57903	=>	10872,
		57904	=>	10874,
		57905	=>	10876,
		57906	=>	10879,
		57907	=>	10881,
		57908	=>	10884,
		57909	=>	10886,
		57910	=>	10888,
		57911	=>	10891,
		57912	=>	10893,
		57913	=>	10895,
		57914	=>	10898,
		57915	=>	10900,
		57916	=>	10902,
		57917	=>	10905,
		57918	=>	10907,
		57919	=>	10909,
		57920	=>	10912,
		57921	=>	10914,
		57922	=>	10916,
		57923	=>	10919,
		57924	=>	10921,
		57925	=>	10923,
		57926	=>	10926,
		57927	=>	10928,
		57928	=>	10930,
		57929	=>	10933,
		57930	=>	10935,
		57931	=>	10937,
		57932	=>	10940,
		57933	=>	10942,
		57934	=>	10944,
		57935	=>	10947,
		57936	=>	10949,
		57937	=>	10951,
		57938	=>	10954,
		57939	=>	10956,
		57940	=>	10958,
		57941	=>	10961,
		57942	=>	10963,
		57943	=>	10965,
		57944	=>	10968,
		57945	=>	10970,
		57946	=>	10973,
		57947	=>	10975,
		57948	=>	10977,
		57949	=>	10980,
		57950	=>	10982,
		57951	=>	10984,
		57952	=>	10987,
		57953	=>	10989,
		57954	=>	10991,
		57955	=>	10994,
		57956	=>	10996,
		57957	=>	10998,
		57958	=>	11001,
		57959	=>	11003,
		57960	=>	11005,
		57961	=>	11008,
		57962	=>	11010,
		57963	=>	11012,
		57964	=>	11015,
		57965	=>	11017,
		57966	=>	11019,
		57967	=>	11022,
		57968	=>	11024,
		57969	=>	11027,
		57970	=>	11029,
		57971	=>	11031,
		57972	=>	11034,
		57973	=>	11036,
		57974	=>	11038,
		57975	=>	11041,
		57976	=>	11043,
		57977	=>	11045,
		57978	=>	11048,
		57979	=>	11050,
		57980	=>	11052,
		57981	=>	11055,
		57982	=>	11057,
		57983	=>	11059,
		57984	=>	11062,
		57985	=>	11064,
		57986	=>	11066,
		57987	=>	11069,
		57988	=>	11071,
		57989	=>	11074,
		57990	=>	11076,
		57991	=>	11078,
		57992	=>	11081,
		57993	=>	11083,
		57994	=>	11085,
		57995	=>	11088,
		57996	=>	11090,
		57997	=>	11092,
		57998	=>	11095,
		57999	=>	11097,
		58000	=>	11099,
		58001	=>	11102,
		58002	=>	11104,
		58003	=>	11107,
		58004	=>	11109,
		58005	=>	11111,
		58006	=>	11114,
		58007	=>	11116,
		58008	=>	11118,
		58009	=>	11121,
		58010	=>	11123,
		58011	=>	11125,
		58012	=>	11128,
		58013	=>	11130,
		58014	=>	11132,
		58015	=>	11135,
		58016	=>	11137,
		58017	=>	11140,
		58018	=>	11142,
		58019	=>	11144,
		58020	=>	11147,
		58021	=>	11149,
		58022	=>	11151,
		58023	=>	11154,
		58024	=>	11156,
		58025	=>	11158,
		58026	=>	11161,
		58027	=>	11163,
		58028	=>	11166,
		58029	=>	11168,
		58030	=>	11170,
		58031	=>	11173,
		58032	=>	11175,
		58033	=>	11177,
		58034	=>	11180,
		58035	=>	11182,
		58036	=>	11184,
		58037	=>	11187,
		58038	=>	11189,
		58039	=>	11192,
		58040	=>	11194,
		58041	=>	11196,
		58042	=>	11199,
		58043	=>	11201,
		58044	=>	11203,
		58045	=>	11206,
		58046	=>	11208,
		58047	=>	11210,
		58048	=>	11213,
		58049	=>	11215,
		58050	=>	11218,
		58051	=>	11220,
		58052	=>	11222,
		58053	=>	11225,
		58054	=>	11227,
		58055	=>	11229,
		58056	=>	11232,
		58057	=>	11234,
		58058	=>	11236,
		58059	=>	11239,
		58060	=>	11241,
		58061	=>	11244,
		58062	=>	11246,
		58063	=>	11248,
		58064	=>	11251,
		58065	=>	11253,
		58066	=>	11255,
		58067	=>	11258,
		58068	=>	11260,
		58069	=>	11263,
		58070	=>	11265,
		58071	=>	11267,
		58072	=>	11270,
		58073	=>	11272,
		58074	=>	11274,
		58075	=>	11277,
		58076	=>	11279,
		58077	=>	11282,
		58078	=>	11284,
		58079	=>	11286,
		58080	=>	11289,
		58081	=>	11291,
		58082	=>	11293,
		58083	=>	11296,
		58084	=>	11298,
		58085	=>	11301,
		58086	=>	11303,
		58087	=>	11305,
		58088	=>	11308,
		58089	=>	11310,
		58090	=>	11312,
		58091	=>	11315,
		58092	=>	11317,
		58093	=>	11319,
		58094	=>	11322,
		58095	=>	11324,
		58096	=>	11327,
		58097	=>	11329,
		58098	=>	11331,
		58099	=>	11334,
		58100	=>	11336,
		58101	=>	11339,
		58102	=>	11341,
		58103	=>	11343,
		58104	=>	11346,
		58105	=>	11348,
		58106	=>	11350,
		58107	=>	11353,
		58108	=>	11355,
		58109	=>	11358,
		58110	=>	11360,
		58111	=>	11362,
		58112	=>	11365,
		58113	=>	11367,
		58114	=>	11369,
		58115	=>	11372,
		58116	=>	11374,
		58117	=>	11377,
		58118	=>	11379,
		58119	=>	11381,
		58120	=>	11384,
		58121	=>	11386,
		58122	=>	11388,
		58123	=>	11391,
		58124	=>	11393,
		58125	=>	11396,
		58126	=>	11398,
		58127	=>	11400,
		58128	=>	11403,
		58129	=>	11405,
		58130	=>	11408,
		58131	=>	11410,
		58132	=>	11412,
		58133	=>	11415,
		58134	=>	11417,
		58135	=>	11419,
		58136	=>	11422,
		58137	=>	11424,
		58138	=>	11427,
		58139	=>	11429,
		58140	=>	11431,
		58141	=>	11434,
		58142	=>	11436,
		58143	=>	11438,
		58144	=>	11441,
		58145	=>	11443,
		58146	=>	11446,
		58147	=>	11448,
		58148	=>	11450,
		58149	=>	11453,
		58150	=>	11455,
		58151	=>	11458,
		58152	=>	11460,
		58153	=>	11462,
		58154	=>	11465,
		58155	=>	11467,
		58156	=>	11470,
		58157	=>	11472,
		58158	=>	11474,
		58159	=>	11477,
		58160	=>	11479,
		58161	=>	11481,
		58162	=>	11484,
		58163	=>	11486,
		58164	=>	11489,
		58165	=>	11491,
		58166	=>	11493,
		58167	=>	11496,
		58168	=>	11498,
		58169	=>	11501,
		58170	=>	11503,
		58171	=>	11505,
		58172	=>	11508,
		58173	=>	11510,
		58174	=>	11513,
		58175	=>	11515,
		58176	=>	11517,
		58177	=>	11520,
		58178	=>	11522,
		58179	=>	11524,
		58180	=>	11527,
		58181	=>	11529,
		58182	=>	11532,
		58183	=>	11534,
		58184	=>	11536,
		58185	=>	11539,
		58186	=>	11541,
		58187	=>	11544,
		58188	=>	11546,
		58189	=>	11548,
		58190	=>	11551,
		58191	=>	11553,
		58192	=>	11556,
		58193	=>	11558,
		58194	=>	11560,
		58195	=>	11563,
		58196	=>	11565,
		58197	=>	11568,
		58198	=>	11570,
		58199	=>	11572,
		58200	=>	11575,
		58201	=>	11577,
		58202	=>	11580,
		58203	=>	11582,
		58204	=>	11584,
		58205	=>	11587,
		58206	=>	11589,
		58207	=>	11592,
		58208	=>	11594,
		58209	=>	11596,
		58210	=>	11599,
		58211	=>	11601,
		58212	=>	11604,
		58213	=>	11606,
		58214	=>	11608,
		58215	=>	11611,
		58216	=>	11613,
		58217	=>	11616,
		58218	=>	11618,
		58219	=>	11620,
		58220	=>	11623,
		58221	=>	11625,
		58222	=>	11628,
		58223	=>	11630,
		58224	=>	11632,
		58225	=>	11635,
		58226	=>	11637,
		58227	=>	11640,
		58228	=>	11642,
		58229	=>	11644,
		58230	=>	11647,
		58231	=>	11649,
		58232	=>	11652,
		58233	=>	11654,
		58234	=>	11656,
		58235	=>	11659,
		58236	=>	11661,
		58237	=>	11664,
		58238	=>	11666,
		58239	=>	11668,
		58240	=>	11671,
		58241	=>	11673,
		58242	=>	11676,
		58243	=>	11678,
		58244	=>	11680,
		58245	=>	11683,
		58246	=>	11685,
		58247	=>	11688,
		58248	=>	11690,
		58249	=>	11692,
		58250	=>	11695,
		58251	=>	11697,
		58252	=>	11700,
		58253	=>	11702,
		58254	=>	11704,
		58255	=>	11707,
		58256	=>	11709,
		58257	=>	11712,
		58258	=>	11714,
		58259	=>	11716,
		58260	=>	11719,
		58261	=>	11721,
		58262	=>	11724,
		58263	=>	11726,
		58264	=>	11728,
		58265	=>	11731,
		58266	=>	11733,
		58267	=>	11736,
		58268	=>	11738,
		58269	=>	11741,
		58270	=>	11743,
		58271	=>	11745,
		58272	=>	11748,
		58273	=>	11750,
		58274	=>	11753,
		58275	=>	11755,
		58276	=>	11757,
		58277	=>	11760,
		58278	=>	11762,
		58279	=>	11765,
		58280	=>	11767,
		58281	=>	11769,
		58282	=>	11772,
		58283	=>	11774,
		58284	=>	11777,
		58285	=>	11779,
		58286	=>	11782,
		58287	=>	11784,
		58288	=>	11786,
		58289	=>	11789,
		58290	=>	11791,
		58291	=>	11794,
		58292	=>	11796,
		58293	=>	11798,
		58294	=>	11801,
		58295	=>	11803,
		58296	=>	11806,
		58297	=>	11808,
		58298	=>	11810,
		58299	=>	11813,
		58300	=>	11815,
		58301	=>	11818,
		58302	=>	11820,
		58303	=>	11823,
		58304	=>	11825,
		58305	=>	11827,
		58306	=>	11830,
		58307	=>	11832,
		58308	=>	11835,
		58309	=>	11837,
		58310	=>	11839,
		58311	=>	11842,
		58312	=>	11844,
		58313	=>	11847,
		58314	=>	11849,
		58315	=>	11852,
		58316	=>	11854,
		58317	=>	11856,
		58318	=>	11859,
		58319	=>	11861,
		58320	=>	11864,
		58321	=>	11866,
		58322	=>	11869,
		58323	=>	11871,
		58324	=>	11873,
		58325	=>	11876,
		58326	=>	11878,
		58327	=>	11881,
		58328	=>	11883,
		58329	=>	11885,
		58330	=>	11888,
		58331	=>	11890,
		58332	=>	11893,
		58333	=>	11895,
		58334	=>	11898,
		58335	=>	11900,
		58336	=>	11902,
		58337	=>	11905,
		58338	=>	11907,
		58339	=>	11910,
		58340	=>	11912,
		58341	=>	11915,
		58342	=>	11917,
		58343	=>	11919,
		58344	=>	11922,
		58345	=>	11924,
		58346	=>	11927,
		58347	=>	11929,
		58348	=>	11931,
		58349	=>	11934,
		58350	=>	11936,
		58351	=>	11939,
		58352	=>	11941,
		58353	=>	11944,
		58354	=>	11946,
		58355	=>	11948,
		58356	=>	11951,
		58357	=>	11953,
		58358	=>	11956,
		58359	=>	11958,
		58360	=>	11961,
		58361	=>	11963,
		58362	=>	11965,
		58363	=>	11968,
		58364	=>	11970,
		58365	=>	11973,
		58366	=>	11975,
		58367	=>	11978,
		58368	=>	11980,
		58369	=>	11982,
		58370	=>	11985,
		58371	=>	11987,
		58372	=>	11990,
		58373	=>	11992,
		58374	=>	11995,
		58375	=>	11997,
		58376	=>	11999,
		58377	=>	12002,
		58378	=>	12004,
		58379	=>	12007,
		58380	=>	12009,
		58381	=>	12012,
		58382	=>	12014,
		58383	=>	12016,
		58384	=>	12019,
		58385	=>	12021,
		58386	=>	12024,
		58387	=>	12026,
		58388	=>	12029,
		58389	=>	12031,
		58390	=>	12033,
		58391	=>	12036,
		58392	=>	12038,
		58393	=>	12041,
		58394	=>	12043,
		58395	=>	12046,
		58396	=>	12048,
		58397	=>	12051,
		58398	=>	12053,
		58399	=>	12055,
		58400	=>	12058,
		58401	=>	12060,
		58402	=>	12063,
		58403	=>	12065,
		58404	=>	12068,
		58405	=>	12070,
		58406	=>	12072,
		58407	=>	12075,
		58408	=>	12077,
		58409	=>	12080,
		58410	=>	12082,
		58411	=>	12085,
		58412	=>	12087,
		58413	=>	12089,
		58414	=>	12092,
		58415	=>	12094,
		58416	=>	12097,
		58417	=>	12099,
		58418	=>	12102,
		58419	=>	12104,
		58420	=>	12107,
		58421	=>	12109,
		58422	=>	12111,
		58423	=>	12114,
		58424	=>	12116,
		58425	=>	12119,
		58426	=>	12121,
		58427	=>	12124,
		58428	=>	12126,
		58429	=>	12129,
		58430	=>	12131,
		58431	=>	12133,
		58432	=>	12136,
		58433	=>	12138,
		58434	=>	12141,
		58435	=>	12143,
		58436	=>	12146,
		58437	=>	12148,
		58438	=>	12150,
		58439	=>	12153,
		58440	=>	12155,
		58441	=>	12158,
		58442	=>	12160,
		58443	=>	12163,
		58444	=>	12165,
		58445	=>	12168,
		58446	=>	12170,
		58447	=>	12172,
		58448	=>	12175,
		58449	=>	12177,
		58450	=>	12180,
		58451	=>	12182,
		58452	=>	12185,
		58453	=>	12187,
		58454	=>	12190,
		58455	=>	12192,
		58456	=>	12194,
		58457	=>	12197,
		58458	=>	12199,
		58459	=>	12202,
		58460	=>	12204,
		58461	=>	12207,
		58462	=>	12209,
		58463	=>	12212,
		58464	=>	12214,
		58465	=>	12216,
		58466	=>	12219,
		58467	=>	12221,
		58468	=>	12224,
		58469	=>	12226,
		58470	=>	12229,
		58471	=>	12231,
		58472	=>	12234,
		58473	=>	12236,
		58474	=>	12239,
		58475	=>	12241,
		58476	=>	12243,
		58477	=>	12246,
		58478	=>	12248,
		58479	=>	12251,
		58480	=>	12253,
		58481	=>	12256,
		58482	=>	12258,
		58483	=>	12261,
		58484	=>	12263,
		58485	=>	12265,
		58486	=>	12268,
		58487	=>	12270,
		58488	=>	12273,
		58489	=>	12275,
		58490	=>	12278,
		58491	=>	12280,
		58492	=>	12283,
		58493	=>	12285,
		58494	=>	12288,
		58495	=>	12290,
		58496	=>	12292,
		58497	=>	12295,
		58498	=>	12297,
		58499	=>	12300,
		58500	=>	12302,
		58501	=>	12305,
		58502	=>	12307,
		58503	=>	12310,
		58504	=>	12312,
		58505	=>	12314,
		58506	=>	12317,
		58507	=>	12319,
		58508	=>	12322,
		58509	=>	12324,
		58510	=>	12327,
		58511	=>	12329,
		58512	=>	12332,
		58513	=>	12334,
		58514	=>	12337,
		58515	=>	12339,
		58516	=>	12342,
		58517	=>	12344,
		58518	=>	12346,
		58519	=>	12349,
		58520	=>	12351,
		58521	=>	12354,
		58522	=>	12356,
		58523	=>	12359,
		58524	=>	12361,
		58525	=>	12364,
		58526	=>	12366,
		58527	=>	12369,
		58528	=>	12371,
		58529	=>	12373,
		58530	=>	12376,
		58531	=>	12378,
		58532	=>	12381,
		58533	=>	12383,
		58534	=>	12386,
		58535	=>	12388,
		58536	=>	12391,
		58537	=>	12393,
		58538	=>	12396,
		58539	=>	12398,
		58540	=>	12401,
		58541	=>	12403,
		58542	=>	12405,
		58543	=>	12408,
		58544	=>	12410,
		58545	=>	12413,
		58546	=>	12415,
		58547	=>	12418,
		58548	=>	12420,
		58549	=>	12423,
		58550	=>	12425,
		58551	=>	12428,
		58552	=>	12430,
		58553	=>	12433,
		58554	=>	12435,
		58555	=>	12437,
		58556	=>	12440,
		58557	=>	12442,
		58558	=>	12445,
		58559	=>	12447,
		58560	=>	12450,
		58561	=>	12452,
		58562	=>	12455,
		58563	=>	12457,
		58564	=>	12460,
		58565	=>	12462,
		58566	=>	12465,
		58567	=>	12467,
		58568	=>	12469,
		58569	=>	12472,
		58570	=>	12474,
		58571	=>	12477,
		58572	=>	12479,
		58573	=>	12482,
		58574	=>	12484,
		58575	=>	12487,
		58576	=>	12489,
		58577	=>	12492,
		58578	=>	12494,
		58579	=>	12497,
		58580	=>	12499,
		58581	=>	12502,
		58582	=>	12504,
		58583	=>	12507,
		58584	=>	12509,
		58585	=>	12511,
		58586	=>	12514,
		58587	=>	12516,
		58588	=>	12519,
		58589	=>	12521,
		58590	=>	12524,
		58591	=>	12526,
		58592	=>	12529,
		58593	=>	12531,
		58594	=>	12534,
		58595	=>	12536,
		58596	=>	12539,
		58597	=>	12541,
		58598	=>	12544,
		58599	=>	12546,
		58600	=>	12549,
		58601	=>	12551,
		58602	=>	12553,
		58603	=>	12556,
		58604	=>	12558,
		58605	=>	12561,
		58606	=>	12563,
		58607	=>	12566,
		58608	=>	12568,
		58609	=>	12571,
		58610	=>	12573,
		58611	=>	12576,
		58612	=>	12578,
		58613	=>	12581,
		58614	=>	12583,
		58615	=>	12586,
		58616	=>	12588,
		58617	=>	12591,
		58618	=>	12593,
		58619	=>	12596,
		58620	=>	12598,
		58621	=>	12600,
		58622	=>	12603,
		58623	=>	12605,
		58624	=>	12608,
		58625	=>	12610,
		58626	=>	12613,
		58627	=>	12615,
		58628	=>	12618,
		58629	=>	12620,
		58630	=>	12623,
		58631	=>	12625,
		58632	=>	12628,
		58633	=>	12630,
		58634	=>	12633,
		58635	=>	12635,
		58636	=>	12638,
		58637	=>	12640,
		58638	=>	12643,
		58639	=>	12645,
		58640	=>	12648,
		58641	=>	12650,
		58642	=>	12653,
		58643	=>	12655,
		58644	=>	12657,
		58645	=>	12660,
		58646	=>	12662,
		58647	=>	12665,
		58648	=>	12667,
		58649	=>	12670,
		58650	=>	12672,
		58651	=>	12675,
		58652	=>	12677,
		58653	=>	12680,
		58654	=>	12682,
		58655	=>	12685,
		58656	=>	12687,
		58657	=>	12690,
		58658	=>	12692,
		58659	=>	12695,
		58660	=>	12697,
		58661	=>	12700,
		58662	=>	12702,
		58663	=>	12705,
		58664	=>	12707,
		58665	=>	12710,
		58666	=>	12712,
		58667	=>	12715,
		58668	=>	12717,
		58669	=>	12720,
		58670	=>	12722,
		58671	=>	12725,
		58672	=>	12727,
		58673	=>	12729,
		58674	=>	12732,
		58675	=>	12734,
		58676	=>	12737,
		58677	=>	12739,
		58678	=>	12742,
		58679	=>	12744,
		58680	=>	12747,
		58681	=>	12749,
		58682	=>	12752,
		58683	=>	12754,
		58684	=>	12757,
		58685	=>	12759,
		58686	=>	12762,
		58687	=>	12764,
		58688	=>	12767,
		58689	=>	12769,
		58690	=>	12772,
		58691	=>	12774,
		58692	=>	12777,
		58693	=>	12779,
		58694	=>	12782,
		58695	=>	12784,
		58696	=>	12787,
		58697	=>	12789,
		58698	=>	12792,
		58699	=>	12794,
		58700	=>	12797,
		58701	=>	12799,
		58702	=>	12802,
		58703	=>	12804,
		58704	=>	12807,
		58705	=>	12809,
		58706	=>	12812,
		58707	=>	12814,
		58708	=>	12817,
		58709	=>	12819,
		58710	=>	12822,
		58711	=>	12824,
		58712	=>	12827,
		58713	=>	12829,
		58714	=>	12832,
		58715	=>	12834,
		58716	=>	12837,
		58717	=>	12839,
		58718	=>	12842,
		58719	=>	12844,
		58720	=>	12847,
		58721	=>	12849,
		58722	=>	12851,
		58723	=>	12854,
		58724	=>	12856,
		58725	=>	12859,
		58726	=>	12861,
		58727	=>	12864,
		58728	=>	12866,
		58729	=>	12869,
		58730	=>	12871,
		58731	=>	12874,
		58732	=>	12876,
		58733	=>	12879,
		58734	=>	12881,
		58735	=>	12884,
		58736	=>	12886,
		58737	=>	12889,
		58738	=>	12891,
		58739	=>	12894,
		58740	=>	12896,
		58741	=>	12899,
		58742	=>	12901,
		58743	=>	12904,
		58744	=>	12906,
		58745	=>	12909,
		58746	=>	12911,
		58747	=>	12914,
		58748	=>	12916,
		58749	=>	12919,
		58750	=>	12921,
		58751	=>	12924,
		58752	=>	12926,
		58753	=>	12929,
		58754	=>	12931,
		58755	=>	12934,
		58756	=>	12936,
		58757	=>	12939,
		58758	=>	12941,
		58759	=>	12944,
		58760	=>	12946,
		58761	=>	12949,
		58762	=>	12951,
		58763	=>	12954,
		58764	=>	12956,
		58765	=>	12959,
		58766	=>	12961,
		58767	=>	12964,
		58768	=>	12966,
		58769	=>	12969,
		58770	=>	12971,
		58771	=>	12974,
		58772	=>	12976,
		58773	=>	12979,
		58774	=>	12981,
		58775	=>	12984,
		58776	=>	12986,
		58777	=>	12989,
		58778	=>	12991,
		58779	=>	12994,
		58780	=>	12996,
		58781	=>	12999,
		58782	=>	13002,
		58783	=>	13004,
		58784	=>	13007,
		58785	=>	13009,
		58786	=>	13012,
		58787	=>	13014,
		58788	=>	13017,
		58789	=>	13019,
		58790	=>	13022,
		58791	=>	13024,
		58792	=>	13027,
		58793	=>	13029,
		58794	=>	13032,
		58795	=>	13034,
		58796	=>	13037,
		58797	=>	13039,
		58798	=>	13042,
		58799	=>	13044,
		58800	=>	13047,
		58801	=>	13049,
		58802	=>	13052,
		58803	=>	13054,
		58804	=>	13057,
		58805	=>	13059,
		58806	=>	13062,
		58807	=>	13064,
		58808	=>	13067,
		58809	=>	13069,
		58810	=>	13072,
		58811	=>	13074,
		58812	=>	13077,
		58813	=>	13079,
		58814	=>	13082,
		58815	=>	13084,
		58816	=>	13087,
		58817	=>	13089,
		58818	=>	13092,
		58819	=>	13094,
		58820	=>	13097,
		58821	=>	13099,
		58822	=>	13102,
		58823	=>	13104,
		58824	=>	13107,
		58825	=>	13109,
		58826	=>	13112,
		58827	=>	13114,
		58828	=>	13117,
		58829	=>	13119,
		58830	=>	13122,
		58831	=>	13124,
		58832	=>	13127,
		58833	=>	13130,
		58834	=>	13132,
		58835	=>	13135,
		58836	=>	13137,
		58837	=>	13140,
		58838	=>	13142,
		58839	=>	13145,
		58840	=>	13147,
		58841	=>	13150,
		58842	=>	13152,
		58843	=>	13155,
		58844	=>	13157,
		58845	=>	13160,
		58846	=>	13162,
		58847	=>	13165,
		58848	=>	13167,
		58849	=>	13170,
		58850	=>	13172,
		58851	=>	13175,
		58852	=>	13177,
		58853	=>	13180,
		58854	=>	13182,
		58855	=>	13185,
		58856	=>	13187,
		58857	=>	13190,
		58858	=>	13192,
		58859	=>	13195,
		58860	=>	13197,
		58861	=>	13200,
		58862	=>	13203,
		58863	=>	13205,
		58864	=>	13208,
		58865	=>	13210,
		58866	=>	13213,
		58867	=>	13215,
		58868	=>	13218,
		58869	=>	13220,
		58870	=>	13223,
		58871	=>	13225,
		58872	=>	13228,
		58873	=>	13230,
		58874	=>	13233,
		58875	=>	13235,
		58876	=>	13238,
		58877	=>	13240,
		58878	=>	13243,
		58879	=>	13245,
		58880	=>	13248,
		58881	=>	13250,
		58882	=>	13253,
		58883	=>	13255,
		58884	=>	13258,
		58885	=>	13261,
		58886	=>	13263,
		58887	=>	13266,
		58888	=>	13268,
		58889	=>	13271,
		58890	=>	13273,
		58891	=>	13276,
		58892	=>	13278,
		58893	=>	13281,
		58894	=>	13283,
		58895	=>	13286,
		58896	=>	13288,
		58897	=>	13291,
		58898	=>	13293,
		58899	=>	13296,
		58900	=>	13298,
		58901	=>	13301,
		58902	=>	13303,
		58903	=>	13306,
		58904	=>	13309,
		58905	=>	13311,
		58906	=>	13314,
		58907	=>	13316,
		58908	=>	13319,
		58909	=>	13321,
		58910	=>	13324,
		58911	=>	13326,
		58912	=>	13329,
		58913	=>	13331,
		58914	=>	13334,
		58915	=>	13336,
		58916	=>	13339,
		58917	=>	13341,
		58918	=>	13344,
		58919	=>	13346,
		58920	=>	13349,
		58921	=>	13352,
		58922	=>	13354,
		58923	=>	13357,
		58924	=>	13359,
		58925	=>	13362,
		58926	=>	13364,
		58927	=>	13367,
		58928	=>	13369,
		58929	=>	13372,
		58930	=>	13374,
		58931	=>	13377,
		58932	=>	13379,
		58933	=>	13382,
		58934	=>	13384,
		58935	=>	13387,
		58936	=>	13390,
		58937	=>	13392,
		58938	=>	13395,
		58939	=>	13397,
		58940	=>	13400,
		58941	=>	13402,
		58942	=>	13405,
		58943	=>	13407,
		58944	=>	13410,
		58945	=>	13412,
		58946	=>	13415,
		58947	=>	13417,
		58948	=>	13420,
		58949	=>	13422,
		58950	=>	13425,
		58951	=>	13428,
		58952	=>	13430,
		58953	=>	13433,
		58954	=>	13435,
		58955	=>	13438,
		58956	=>	13440,
		58957	=>	13443,
		58958	=>	13445,
		58959	=>	13448,
		58960	=>	13450,
		58961	=>	13453,
		58962	=>	13455,
		58963	=>	13458,
		58964	=>	13461,
		58965	=>	13463,
		58966	=>	13466,
		58967	=>	13468,
		58968	=>	13471,
		58969	=>	13473,
		58970	=>	13476,
		58971	=>	13478,
		58972	=>	13481,
		58973	=>	13483,
		58974	=>	13486,
		58975	=>	13488,
		58976	=>	13491,
		58977	=>	13494,
		58978	=>	13496,
		58979	=>	13499,
		58980	=>	13501,
		58981	=>	13504,
		58982	=>	13506,
		58983	=>	13509,
		58984	=>	13511,
		58985	=>	13514,
		58986	=>	13516,
		58987	=>	13519,
		58988	=>	13521,
		58989	=>	13524,
		58990	=>	13527,
		58991	=>	13529,
		58992	=>	13532,
		58993	=>	13534,
		58994	=>	13537,
		58995	=>	13539,
		58996	=>	13542,
		58997	=>	13544,
		58998	=>	13547,
		58999	=>	13549,
		59000	=>	13552,
		59001	=>	13555,
		59002	=>	13557,
		59003	=>	13560,
		59004	=>	13562,
		59005	=>	13565,
		59006	=>	13567,
		59007	=>	13570,
		59008	=>	13572,
		59009	=>	13575,
		59010	=>	13577,
		59011	=>	13580,
		59012	=>	13583,
		59013	=>	13585,
		59014	=>	13588,
		59015	=>	13590,
		59016	=>	13593,
		59017	=>	13595,
		59018	=>	13598,
		59019	=>	13600,
		59020	=>	13603,
		59021	=>	13605,
		59022	=>	13608,
		59023	=>	13611,
		59024	=>	13613,
		59025	=>	13616,
		59026	=>	13618,
		59027	=>	13621,
		59028	=>	13623,
		59029	=>	13626,
		59030	=>	13628,
		59031	=>	13631,
		59032	=>	13634,
		59033	=>	13636,
		59034	=>	13639,
		59035	=>	13641,
		59036	=>	13644,
		59037	=>	13646,
		59038	=>	13649,
		59039	=>	13651,
		59040	=>	13654,
		59041	=>	13656,
		59042	=>	13659,
		59043	=>	13662,
		59044	=>	13664,
		59045	=>	13667,
		59046	=>	13669,
		59047	=>	13672,
		59048	=>	13674,
		59049	=>	13677,
		59050	=>	13679,
		59051	=>	13682,
		59052	=>	13685,
		59053	=>	13687,
		59054	=>	13690,
		59055	=>	13692,
		59056	=>	13695,
		59057	=>	13697,
		59058	=>	13700,
		59059	=>	13702,
		59060	=>	13705,
		59061	=>	13708,
		59062	=>	13710,
		59063	=>	13713,
		59064	=>	13715,
		59065	=>	13718,
		59066	=>	13720,
		59067	=>	13723,
		59068	=>	13725,
		59069	=>	13728,
		59070	=>	13731,
		59071	=>	13733,
		59072	=>	13736,
		59073	=>	13738,
		59074	=>	13741,
		59075	=>	13743,
		59076	=>	13746,
		59077	=>	13748,
		59078	=>	13751,
		59079	=>	13754,
		59080	=>	13756,
		59081	=>	13759,
		59082	=>	13761,
		59083	=>	13764,
		59084	=>	13766,
		59085	=>	13769,
		59086	=>	13771,
		59087	=>	13774,
		59088	=>	13777,
		59089	=>	13779,
		59090	=>	13782,
		59091	=>	13784,
		59092	=>	13787,
		59093	=>	13789,
		59094	=>	13792,
		59095	=>	13795,
		59096	=>	13797,
		59097	=>	13800,
		59098	=>	13802,
		59099	=>	13805,
		59100	=>	13807,
		59101	=>	13810,
		59102	=>	13812,
		59103	=>	13815,
		59104	=>	13818,
		59105	=>	13820,
		59106	=>	13823,
		59107	=>	13825,
		59108	=>	13828,
		59109	=>	13830,
		59110	=>	13833,
		59111	=>	13836,
		59112	=>	13838,
		59113	=>	13841,
		59114	=>	13843,
		59115	=>	13846,
		59116	=>	13848,
		59117	=>	13851,
		59118	=>	13854,
		59119	=>	13856,
		59120	=>	13859,
		59121	=>	13861,
		59122	=>	13864,
		59123	=>	13866,
		59124	=>	13869,
		59125	=>	13871,
		59126	=>	13874,
		59127	=>	13877,
		59128	=>	13879,
		59129	=>	13882,
		59130	=>	13884,
		59131	=>	13887,
		59132	=>	13889,
		59133	=>	13892,
		59134	=>	13895,
		59135	=>	13897,
		59136	=>	13900,
		59137	=>	13902,
		59138	=>	13905,
		59139	=>	13907,
		59140	=>	13910,
		59141	=>	13913,
		59142	=>	13915,
		59143	=>	13918,
		59144	=>	13920,
		59145	=>	13923,
		59146	=>	13925,
		59147	=>	13928,
		59148	=>	13931,
		59149	=>	13933,
		59150	=>	13936,
		59151	=>	13938,
		59152	=>	13941,
		59153	=>	13943,
		59154	=>	13946,
		59155	=>	13949,
		59156	=>	13951,
		59157	=>	13954,
		59158	=>	13956,
		59159	=>	13959,
		59160	=>	13961,
		59161	=>	13964,
		59162	=>	13967,
		59163	=>	13969,
		59164	=>	13972,
		59165	=>	13974,
		59166	=>	13977,
		59167	=>	13979,
		59168	=>	13982,
		59169	=>	13985,
		59170	=>	13987,
		59171	=>	13990,
		59172	=>	13992,
		59173	=>	13995,
		59174	=>	13997,
		59175	=>	14000,
		59176	=>	14003,
		59177	=>	14005,
		59178	=>	14008,
		59179	=>	14010,
		59180	=>	14013,
		59181	=>	14015,
		59182	=>	14018,
		59183	=>	14021,
		59184	=>	14023,
		59185	=>	14026,
		59186	=>	14028,
		59187	=>	14031,
		59188	=>	14033,
		59189	=>	14036,
		59190	=>	14039,
		59191	=>	14041,
		59192	=>	14044,
		59193	=>	14046,
		59194	=>	14049,
		59195	=>	14052,
		59196	=>	14054,
		59197	=>	14057,
		59198	=>	14059,
		59199	=>	14062,
		59200	=>	14064,
		59201	=>	14067,
		59202	=>	14070,
		59203	=>	14072,
		59204	=>	14075,
		59205	=>	14077,
		59206	=>	14080,
		59207	=>	14083,
		59208	=>	14085,
		59209	=>	14088,
		59210	=>	14090,
		59211	=>	14093,
		59212	=>	14095,
		59213	=>	14098,
		59214	=>	14101,
		59215	=>	14103,
		59216	=>	14106,
		59217	=>	14108,
		59218	=>	14111,
		59219	=>	14113,
		59220	=>	14116,
		59221	=>	14119,
		59222	=>	14121,
		59223	=>	14124,
		59224	=>	14126,
		59225	=>	14129,
		59226	=>	14132,
		59227	=>	14134,
		59228	=>	14137,
		59229	=>	14139,
		59230	=>	14142,
		59231	=>	14144,
		59232	=>	14147,
		59233	=>	14150,
		59234	=>	14152,
		59235	=>	14155,
		59236	=>	14157,
		59237	=>	14160,
		59238	=>	14163,
		59239	=>	14165,
		59240	=>	14168,
		59241	=>	14170,
		59242	=>	14173,
		59243	=>	14176,
		59244	=>	14178,
		59245	=>	14181,
		59246	=>	14183,
		59247	=>	14186,
		59248	=>	14188,
		59249	=>	14191,
		59250	=>	14194,
		59251	=>	14196,
		59252	=>	14199,
		59253	=>	14201,
		59254	=>	14204,
		59255	=>	14207,
		59256	=>	14209,
		59257	=>	14212,
		59258	=>	14214,
		59259	=>	14217,
		59260	=>	14220,
		59261	=>	14222,
		59262	=>	14225,
		59263	=>	14227,
		59264	=>	14230,
		59265	=>	14232,
		59266	=>	14235,
		59267	=>	14238,
		59268	=>	14240,
		59269	=>	14243,
		59270	=>	14245,
		59271	=>	14248,
		59272	=>	14251,
		59273	=>	14253,
		59274	=>	14256,
		59275	=>	14258,
		59276	=>	14261,
		59277	=>	14264,
		59278	=>	14266,
		59279	=>	14269,
		59280	=>	14271,
		59281	=>	14274,
		59282	=>	14277,
		59283	=>	14279,
		59284	=>	14282,
		59285	=>	14284,
		59286	=>	14287,
		59287	=>	14290,
		59288	=>	14292,
		59289	=>	14295,
		59290	=>	14297,
		59291	=>	14300,
		59292	=>	14302,
		59293	=>	14305,
		59294	=>	14308,
		59295	=>	14310,
		59296	=>	14313,
		59297	=>	14315,
		59298	=>	14318,
		59299	=>	14321,
		59300	=>	14323,
		59301	=>	14326,
		59302	=>	14328,
		59303	=>	14331,
		59304	=>	14334,
		59305	=>	14336,
		59306	=>	14339,
		59307	=>	14341,
		59308	=>	14344,
		59309	=>	14347,
		59310	=>	14349,
		59311	=>	14352,
		59312	=>	14354,
		59313	=>	14357,
		59314	=>	14360,
		59315	=>	14362,
		59316	=>	14365,
		59317	=>	14367,
		59318	=>	14370,
		59319	=>	14373,
		59320	=>	14375,
		59321	=>	14378,
		59322	=>	14380,
		59323	=>	14383,
		59324	=>	14386,
		59325	=>	14388,
		59326	=>	14391,
		59327	=>	14393,
		59328	=>	14396,
		59329	=>	14399,
		59330	=>	14401,
		59331	=>	14404,
		59332	=>	14406,
		59333	=>	14409,
		59334	=>	14412,
		59335	=>	14414,
		59336	=>	14417,
		59337	=>	14419,
		59338	=>	14422,
		59339	=>	14425,
		59340	=>	14427,
		59341	=>	14430,
		59342	=>	14432,
		59343	=>	14435,
		59344	=>	14438,
		59345	=>	14440,
		59346	=>	14443,
		59347	=>	14445,
		59348	=>	14448,
		59349	=>	14451,
		59350	=>	14453,
		59351	=>	14456,
		59352	=>	14459,
		59353	=>	14461,
		59354	=>	14464,
		59355	=>	14466,
		59356	=>	14469,
		59357	=>	14472,
		59358	=>	14474,
		59359	=>	14477,
		59360	=>	14479,
		59361	=>	14482,
		59362	=>	14485,
		59363	=>	14487,
		59364	=>	14490,
		59365	=>	14492,
		59366	=>	14495,
		59367	=>	14498,
		59368	=>	14500,
		59369	=>	14503,
		59370	=>	14505,
		59371	=>	14508,
		59372	=>	14511,
		59373	=>	14513,
		59374	=>	14516,
		59375	=>	14518,
		59376	=>	14521,
		59377	=>	14524,
		59378	=>	14526,
		59379	=>	14529,
		59380	=>	14532,
		59381	=>	14534,
		59382	=>	14537,
		59383	=>	14539,
		59384	=>	14542,
		59385	=>	14545,
		59386	=>	14547,
		59387	=>	14550,
		59388	=>	14552,
		59389	=>	14555,
		59390	=>	14558,
		59391	=>	14560,
		59392	=>	14563,
		59393	=>	14565,
		59394	=>	14568,
		59395	=>	14571,
		59396	=>	14573,
		59397	=>	14576,
		59398	=>	14579,
		59399	=>	14581,
		59400	=>	14584,
		59401	=>	14586,
		59402	=>	14589,
		59403	=>	14592,
		59404	=>	14594,
		59405	=>	14597,
		59406	=>	14599,
		59407	=>	14602,
		59408	=>	14605,
		59409	=>	14607,
		59410	=>	14610,
		59411	=>	14613,
		59412	=>	14615,
		59413	=>	14618,
		59414	=>	14620,
		59415	=>	14623,
		59416	=>	14626,
		59417	=>	14628,
		59418	=>	14631,
		59419	=>	14633,
		59420	=>	14636,
		59421	=>	14639,
		59422	=>	14641,
		59423	=>	14644,
		59424	=>	14647,
		59425	=>	14649,
		59426	=>	14652,
		59427	=>	14654,
		59428	=>	14657,
		59429	=>	14660,
		59430	=>	14662,
		59431	=>	14665,
		59432	=>	14667,
		59433	=>	14670,
		59434	=>	14673,
		59435	=>	14675,
		59436	=>	14678,
		59437	=>	14681,
		59438	=>	14683,
		59439	=>	14686,
		59440	=>	14688,
		59441	=>	14691,
		59442	=>	14694,
		59443	=>	14696,
		59444	=>	14699,
		59445	=>	14702,
		59446	=>	14704,
		59447	=>	14707,
		59448	=>	14709,
		59449	=>	14712,
		59450	=>	14715,
		59451	=>	14717,
		59452	=>	14720,
		59453	=>	14723,
		59454	=>	14725,
		59455	=>	14728,
		59456	=>	14730,
		59457	=>	14733,
		59458	=>	14736,
		59459	=>	14738,
		59460	=>	14741,
		59461	=>	14743,
		59462	=>	14746,
		59463	=>	14749,
		59464	=>	14751,
		59465	=>	14754,
		59466	=>	14757,
		59467	=>	14759,
		59468	=>	14762,
		59469	=>	14764,
		59470	=>	14767,
		59471	=>	14770,
		59472	=>	14772,
		59473	=>	14775,
		59474	=>	14778,
		59475	=>	14780,
		59476	=>	14783,
		59477	=>	14785,
		59478	=>	14788,
		59479	=>	14791,
		59480	=>	14793,
		59481	=>	14796,
		59482	=>	14799,
		59483	=>	14801,
		59484	=>	14804,
		59485	=>	14806,
		59486	=>	14809,
		59487	=>	14812,
		59488	=>	14814,
		59489	=>	14817,
		59490	=>	14820,
		59491	=>	14822,
		59492	=>	14825,
		59493	=>	14828,
		59494	=>	14830,
		59495	=>	14833,
		59496	=>	14835,
		59497	=>	14838,
		59498	=>	14841,
		59499	=>	14843,
		59500	=>	14846,
		59501	=>	14849,
		59502	=>	14851,
		59503	=>	14854,
		59504	=>	14856,
		59505	=>	14859,
		59506	=>	14862,
		59507	=>	14864,
		59508	=>	14867,
		59509	=>	14870,
		59510	=>	14872,
		59511	=>	14875,
		59512	=>	14878,
		59513	=>	14880,
		59514	=>	14883,
		59515	=>	14885,
		59516	=>	14888,
		59517	=>	14891,
		59518	=>	14893,
		59519	=>	14896,
		59520	=>	14899,
		59521	=>	14901,
		59522	=>	14904,
		59523	=>	14906,
		59524	=>	14909,
		59525	=>	14912,
		59526	=>	14914,
		59527	=>	14917,
		59528	=>	14920,
		59529	=>	14922,
		59530	=>	14925,
		59531	=>	14928,
		59532	=>	14930,
		59533	=>	14933,
		59534	=>	14935,
		59535	=>	14938,
		59536	=>	14941,
		59537	=>	14943,
		59538	=>	14946,
		59539	=>	14949,
		59540	=>	14951,
		59541	=>	14954,
		59542	=>	14957,
		59543	=>	14959,
		59544	=>	14962,
		59545	=>	14964,
		59546	=>	14967,
		59547	=>	14970,
		59548	=>	14972,
		59549	=>	14975,
		59550	=>	14978,
		59551	=>	14980,
		59552	=>	14983,
		59553	=>	14986,
		59554	=>	14988,
		59555	=>	14991,
		59556	=>	14993,
		59557	=>	14996,
		59558	=>	14999,
		59559	=>	15001,
		59560	=>	15004,
		59561	=>	15007,
		59562	=>	15009,
		59563	=>	15012,
		59564	=>	15015,
		59565	=>	15017,
		59566	=>	15020,
		59567	=>	15023,
		59568	=>	15025,
		59569	=>	15028,
		59570	=>	15030,
		59571	=>	15033,
		59572	=>	15036,
		59573	=>	15038,
		59574	=>	15041,
		59575	=>	15044,
		59576	=>	15046,
		59577	=>	15049,
		59578	=>	15052,
		59579	=>	15054,
		59580	=>	15057,
		59581	=>	15060,
		59582	=>	15062,
		59583	=>	15065,
		59584	=>	15067,
		59585	=>	15070,
		59586	=>	15073,
		59587	=>	15075,
		59588	=>	15078,
		59589	=>	15081,
		59590	=>	15083,
		59591	=>	15086,
		59592	=>	15089,
		59593	=>	15091,
		59594	=>	15094,
		59595	=>	15097,
		59596	=>	15099,
		59597	=>	15102,
		59598	=>	15104,
		59599	=>	15107,
		59600	=>	15110,
		59601	=>	15112,
		59602	=>	15115,
		59603	=>	15118,
		59604	=>	15120,
		59605	=>	15123,
		59606	=>	15126,
		59607	=>	15128,
		59608	=>	15131,
		59609	=>	15134,
		59610	=>	15136,
		59611	=>	15139,
		59612	=>	15142,
		59613	=>	15144,
		59614	=>	15147,
		59615	=>	15149,
		59616	=>	15152,
		59617	=>	15155,
		59618	=>	15157,
		59619	=>	15160,
		59620	=>	15163,
		59621	=>	15165,
		59622	=>	15168,
		59623	=>	15171,
		59624	=>	15173,
		59625	=>	15176,
		59626	=>	15179,
		59627	=>	15181,
		59628	=>	15184,
		59629	=>	15187,
		59630	=>	15189,
		59631	=>	15192,
		59632	=>	15195,
		59633	=>	15197,
		59634	=>	15200,
		59635	=>	15202,
		59636	=>	15205,
		59637	=>	15208,
		59638	=>	15210,
		59639	=>	15213,
		59640	=>	15216,
		59641	=>	15218,
		59642	=>	15221,
		59643	=>	15224,
		59644	=>	15226,
		59645	=>	15229,
		59646	=>	15232,
		59647	=>	15234,
		59648	=>	15237,
		59649	=>	15240,
		59650	=>	15242,
		59651	=>	15245,
		59652	=>	15248,
		59653	=>	15250,
		59654	=>	15253,
		59655	=>	15256,
		59656	=>	15258,
		59657	=>	15261,
		59658	=>	15264,
		59659	=>	15266,
		59660	=>	15269,
		59661	=>	15271,
		59662	=>	15274,
		59663	=>	15277,
		59664	=>	15279,
		59665	=>	15282,
		59666	=>	15285,
		59667	=>	15287,
		59668	=>	15290,
		59669	=>	15293,
		59670	=>	15295,
		59671	=>	15298,
		59672	=>	15301,
		59673	=>	15303,
		59674	=>	15306,
		59675	=>	15309,
		59676	=>	15311,
		59677	=>	15314,
		59678	=>	15317,
		59679	=>	15319,
		59680	=>	15322,
		59681	=>	15325,
		59682	=>	15327,
		59683	=>	15330,
		59684	=>	15333,
		59685	=>	15335,
		59686	=>	15338,
		59687	=>	15341,
		59688	=>	15343,
		59689	=>	15346,
		59690	=>	15349,
		59691	=>	15351,
		59692	=>	15354,
		59693	=>	15357,
		59694	=>	15359,
		59695	=>	15362,
		59696	=>	15365,
		59697	=>	15367,
		59698	=>	15370,
		59699	=>	15373,
		59700	=>	15375,
		59701	=>	15378,
		59702	=>	15381,
		59703	=>	15383,
		59704	=>	15386,
		59705	=>	15389,
		59706	=>	15391,
		59707	=>	15394,
		59708	=>	15397,
		59709	=>	15399,
		59710	=>	15402,
		59711	=>	15404,
		59712	=>	15407,
		59713	=>	15410,
		59714	=>	15412,
		59715	=>	15415,
		59716	=>	15418,
		59717	=>	15420,
		59718	=>	15423,
		59719	=>	15426,
		59720	=>	15428,
		59721	=>	15431,
		59722	=>	15434,
		59723	=>	15436,
		59724	=>	15439,
		59725	=>	15442,
		59726	=>	15444,
		59727	=>	15447,
		59728	=>	15450,
		59729	=>	15452,
		59730	=>	15455,
		59731	=>	15458,
		59732	=>	15460,
		59733	=>	15463,
		59734	=>	15466,
		59735	=>	15468,
		59736	=>	15471,
		59737	=>	15474,
		59738	=>	15476,
		59739	=>	15479,
		59740	=>	15482,
		59741	=>	15484,
		59742	=>	15487,
		59743	=>	15490,
		59744	=>	15493,
		59745	=>	15495,
		59746	=>	15498,
		59747	=>	15501,
		59748	=>	15503,
		59749	=>	15506,
		59750	=>	15509,
		59751	=>	15511,
		59752	=>	15514,
		59753	=>	15517,
		59754	=>	15519,
		59755	=>	15522,
		59756	=>	15525,
		59757	=>	15527,
		59758	=>	15530,
		59759	=>	15533,
		59760	=>	15535,
		59761	=>	15538,
		59762	=>	15541,
		59763	=>	15543,
		59764	=>	15546,
		59765	=>	15549,
		59766	=>	15551,
		59767	=>	15554,
		59768	=>	15557,
		59769	=>	15559,
		59770	=>	15562,
		59771	=>	15565,
		59772	=>	15567,
		59773	=>	15570,
		59774	=>	15573,
		59775	=>	15575,
		59776	=>	15578,
		59777	=>	15581,
		59778	=>	15583,
		59779	=>	15586,
		59780	=>	15589,
		59781	=>	15591,
		59782	=>	15594,
		59783	=>	15597,
		59784	=>	15599,
		59785	=>	15602,
		59786	=>	15605,
		59787	=>	15607,
		59788	=>	15610,
		59789	=>	15613,
		59790	=>	15615,
		59791	=>	15618,
		59792	=>	15621,
		59793	=>	15623,
		59794	=>	15626,
		59795	=>	15629,
		59796	=>	15632,
		59797	=>	15634,
		59798	=>	15637,
		59799	=>	15640,
		59800	=>	15642,
		59801	=>	15645,
		59802	=>	15648,
		59803	=>	15650,
		59804	=>	15653,
		59805	=>	15656,
		59806	=>	15658,
		59807	=>	15661,
		59808	=>	15664,
		59809	=>	15666,
		59810	=>	15669,
		59811	=>	15672,
		59812	=>	15674,
		59813	=>	15677,
		59814	=>	15680,
		59815	=>	15682,
		59816	=>	15685,
		59817	=>	15688,
		59818	=>	15690,
		59819	=>	15693,
		59820	=>	15696,
		59821	=>	15699,
		59822	=>	15701,
		59823	=>	15704,
		59824	=>	15707,
		59825	=>	15709,
		59826	=>	15712,
		59827	=>	15715,
		59828	=>	15717,
		59829	=>	15720,
		59830	=>	15723,
		59831	=>	15725,
		59832	=>	15728,
		59833	=>	15731,
		59834	=>	15733,
		59835	=>	15736,
		59836	=>	15739,
		59837	=>	15741,
		59838	=>	15744,
		59839	=>	15747,
		59840	=>	15750,
		59841	=>	15752,
		59842	=>	15755,
		59843	=>	15758,
		59844	=>	15760,
		59845	=>	15763,
		59846	=>	15766,
		59847	=>	15768,
		59848	=>	15771,
		59849	=>	15774,
		59850	=>	15776,
		59851	=>	15779,
		59852	=>	15782,
		59853	=>	15784,
		59854	=>	15787,
		59855	=>	15790,
		59856	=>	15792,
		59857	=>	15795,
		59858	=>	15798,
		59859	=>	15801,
		59860	=>	15803,
		59861	=>	15806,
		59862	=>	15809,
		59863	=>	15811,
		59864	=>	15814,
		59865	=>	15817,
		59866	=>	15819,
		59867	=>	15822,
		59868	=>	15825,
		59869	=>	15827,
		59870	=>	15830,
		59871	=>	15833,
		59872	=>	15835,
		59873	=>	15838,
		59874	=>	15841,
		59875	=>	15844,
		59876	=>	15846,
		59877	=>	15849,
		59878	=>	15852,
		59879	=>	15854,
		59880	=>	15857,
		59881	=>	15860,
		59882	=>	15862,
		59883	=>	15865,
		59884	=>	15868,
		59885	=>	15870,
		59886	=>	15873,
		59887	=>	15876,
		59888	=>	15879,
		59889	=>	15881,
		59890	=>	15884,
		59891	=>	15887,
		59892	=>	15889,
		59893	=>	15892,
		59894	=>	15895,
		59895	=>	15897,
		59896	=>	15900,
		59897	=>	15903,
		59898	=>	15905,
		59899	=>	15908,
		59900	=>	15911,
		59901	=>	15914,
		59902	=>	15916,
		59903	=>	15919,
		59904	=>	15922,
		59905	=>	15924,
		59906	=>	15927,
		59907	=>	15930,
		59908	=>	15932,
		59909	=>	15935,
		59910	=>	15938,
		59911	=>	15941,
		59912	=>	15943,
		59913	=>	15946,
		59914	=>	15949,
		59915	=>	15951,
		59916	=>	15954,
		59917	=>	15957,
		59918	=>	15959,
		59919	=>	15962,
		59920	=>	15965,
		59921	=>	15967,
		59922	=>	15970,
		59923	=>	15973,
		59924	=>	15976,
		59925	=>	15978,
		59926	=>	15981,
		59927	=>	15984,
		59928	=>	15986,
		59929	=>	15989,
		59930	=>	15992,
		59931	=>	15994,
		59932	=>	15997,
		59933	=>	16000,
		59934	=>	16003,
		59935	=>	16005,
		59936	=>	16008,
		59937	=>	16011,
		59938	=>	16013,
		59939	=>	16016,
		59940	=>	16019,
		59941	=>	16021,
		59942	=>	16024,
		59943	=>	16027,
		59944	=>	16030,
		59945	=>	16032,
		59946	=>	16035,
		59947	=>	16038,
		59948	=>	16040,
		59949	=>	16043,
		59950	=>	16046,
		59951	=>	16048,
		59952	=>	16051,
		59953	=>	16054,
		59954	=>	16057,
		59955	=>	16059,
		59956	=>	16062,
		59957	=>	16065,
		59958	=>	16067,
		59959	=>	16070,
		59960	=>	16073,
		59961	=>	16075,
		59962	=>	16078,
		59963	=>	16081,
		59964	=>	16084,
		59965	=>	16086,
		59966	=>	16089,
		59967	=>	16092,
		59968	=>	16094,
		59969	=>	16097,
		59970	=>	16100,
		59971	=>	16103,
		59972	=>	16105,
		59973	=>	16108,
		59974	=>	16111,
		59975	=>	16113,
		59976	=>	16116,
		59977	=>	16119,
		59978	=>	16121,
		59979	=>	16124,
		59980	=>	16127,
		59981	=>	16130,
		59982	=>	16132,
		59983	=>	16135,
		59984	=>	16138,
		59985	=>	16140,
		59986	=>	16143,
		59987	=>	16146,
		59988	=>	16149,
		59989	=>	16151,
		59990	=>	16154,
		59991	=>	16157,
		59992	=>	16159,
		59993	=>	16162,
		59994	=>	16165,
		59995	=>	16167,
		59996	=>	16170,
		59997	=>	16173,
		59998	=>	16176,
		59999	=>	16178,
		60000	=>	16181,
		60001	=>	16184,
		60002	=>	16186,
		60003	=>	16189,
		60004	=>	16192,
		60005	=>	16195,
		60006	=>	16197,
		60007	=>	16200,
		60008	=>	16203,
		60009	=>	16205,
		60010	=>	16208,
		60011	=>	16211,
		60012	=>	16214,
		60013	=>	16216,
		60014	=>	16219,
		60015	=>	16222,
		60016	=>	16224,
		60017	=>	16227,
		60018	=>	16230,
		60019	=>	16233,
		60020	=>	16235,
		60021	=>	16238,
		60022	=>	16241,
		60023	=>	16243,
		60024	=>	16246,
		60025	=>	16249,
		60026	=>	16252,
		60027	=>	16254,
		60028	=>	16257,
		60029	=>	16260,
		60030	=>	16262,
		60031	=>	16265,
		60032	=>	16268,
		60033	=>	16271,
		60034	=>	16273,
		60035	=>	16276,
		60036	=>	16279,
		60037	=>	16281,
		60038	=>	16284,
		60039	=>	16287,
		60040	=>	16290,
		60041	=>	16292,
		60042	=>	16295,
		60043	=>	16298,
		60044	=>	16300,
		60045	=>	16303,
		60046	=>	16306,
		60047	=>	16309,
		60048	=>	16311,
		60049	=>	16314,
		60050	=>	16317,
		60051	=>	16319,
		60052	=>	16322,
		60053	=>	16325,
		60054	=>	16328,
		60055	=>	16330,
		60056	=>	16333,
		60057	=>	16336,
		60058	=>	16338,
		60059	=>	16341,
		60060	=>	16344,
		60061	=>	16347,
		60062	=>	16349,
		60063	=>	16352,
		60064	=>	16355,
		60065	=>	16357,
		60066	=>	16360,
		60067	=>	16363,
		60068	=>	16366,
		60069	=>	16368,
		60070	=>	16371,
		60071	=>	16374,
		60072	=>	16376,
		60073	=>	16379,
		60074	=>	16382,
		60075	=>	16385,
		60076	=>	16387,
		60077	=>	16390,
		60078	=>	16393,
		60079	=>	16396,
		60080	=>	16398,
		60081	=>	16401,
		60082	=>	16404,
		60083	=>	16406,
		60084	=>	16409,
		60085	=>	16412,
		60086	=>	16415,
		60087	=>	16417,
		60088	=>	16420,
		60089	=>	16423,
		60090	=>	16425,
		60091	=>	16428,
		60092	=>	16431,
		60093	=>	16434,
		60094	=>	16436,
		60095	=>	16439,
		60096	=>	16442,
		60097	=>	16445,
		60098	=>	16447,
		60099	=>	16450,
		60100	=>	16453,
		60101	=>	16455,
		60102	=>	16458,
		60103	=>	16461,
		60104	=>	16464,
		60105	=>	16466,
		60106	=>	16469,
		60107	=>	16472,
		60108	=>	16475,
		60109	=>	16477,
		60110	=>	16480,
		60111	=>	16483,
		60112	=>	16485,
		60113	=>	16488,
		60114	=>	16491,
		60115	=>	16494,
		60116	=>	16496,
		60117	=>	16499,
		60118	=>	16502,
		60119	=>	16505,
		60120	=>	16507,
		60121	=>	16510,
		60122	=>	16513,
		60123	=>	16515,
		60124	=>	16518,
		60125	=>	16521,
		60126	=>	16524,
		60127	=>	16526,
		60128	=>	16529,
		60129	=>	16532,
		60130	=>	16535,
		60131	=>	16537,
		60132	=>	16540,
		60133	=>	16543,
		60134	=>	16545,
		60135	=>	16548,
		60136	=>	16551,
		60137	=>	16554,
		60138	=>	16556,
		60139	=>	16559,
		60140	=>	16562,
		60141	=>	16565,
		60142	=>	16567,
		60143	=>	16570,
		60144	=>	16573,
		60145	=>	16575,
		60146	=>	16578,
		60147	=>	16581,
		60148	=>	16584,
		60149	=>	16586,
		60150	=>	16589,
		60151	=>	16592,
		60152	=>	16595,
		60153	=>	16597,
		60154	=>	16600,
		60155	=>	16603,
		60156	=>	16606,
		60157	=>	16608,
		60158	=>	16611,
		60159	=>	16614,
		60160	=>	16616,
		60161	=>	16619,
		60162	=>	16622,
		60163	=>	16625,
		60164	=>	16627,
		60165	=>	16630,
		60166	=>	16633,
		60167	=>	16636,
		60168	=>	16638,
		60169	=>	16641,
		60170	=>	16644,
		60171	=>	16647,
		60172	=>	16649,
		60173	=>	16652,
		60174	=>	16655,
		60175	=>	16657,
		60176	=>	16660,
		60177	=>	16663,
		60178	=>	16666,
		60179	=>	16668,
		60180	=>	16671,
		60181	=>	16674,
		60182	=>	16677,
		60183	=>	16679,
		60184	=>	16682,
		60185	=>	16685,
		60186	=>	16688,
		60187	=>	16690,
		60188	=>	16693,
		60189	=>	16696,
		60190	=>	16699,
		60191	=>	16701,
		60192	=>	16704,
		60193	=>	16707,
		60194	=>	16709,
		60195	=>	16712,
		60196	=>	16715,
		60197	=>	16718,
		60198	=>	16720,
		60199	=>	16723,
		60200	=>	16726,
		60201	=>	16729,
		60202	=>	16731,
		60203	=>	16734,
		60204	=>	16737,
		60205	=>	16740,
		60206	=>	16742,
		60207	=>	16745,
		60208	=>	16748,
		60209	=>	16751,
		60210	=>	16753,
		60211	=>	16756,
		60212	=>	16759,
		60213	=>	16762,
		60214	=>	16764,
		60215	=>	16767,
		60216	=>	16770,
		60217	=>	16773,
		60218	=>	16775,
		60219	=>	16778,
		60220	=>	16781,
		60221	=>	16783,
		60222	=>	16786,
		60223	=>	16789,
		60224	=>	16792,
		60225	=>	16794,
		60226	=>	16797,
		60227	=>	16800,
		60228	=>	16803,
		60229	=>	16805,
		60230	=>	16808,
		60231	=>	16811,
		60232	=>	16814,
		60233	=>	16816,
		60234	=>	16819,
		60235	=>	16822,
		60236	=>	16825,
		60237	=>	16827,
		60238	=>	16830,
		60239	=>	16833,
		60240	=>	16836,
		60241	=>	16838,
		60242	=>	16841,
		60243	=>	16844,
		60244	=>	16847,
		60245	=>	16849,
		60246	=>	16852,
		60247	=>	16855,
		60248	=>	16858,
		60249	=>	16860,
		60250	=>	16863,
		60251	=>	16866,
		60252	=>	16869,
		60253	=>	16871,
		60254	=>	16874,
		60255	=>	16877,
		60256	=>	16880,
		60257	=>	16882,
		60258	=>	16885,
		60259	=>	16888,
		60260	=>	16891,
		60261	=>	16893,
		60262	=>	16896,
		60263	=>	16899,
		60264	=>	16902,
		60265	=>	16904,
		60266	=>	16907,
		60267	=>	16910,
		60268	=>	16913,
		60269	=>	16915,
		60270	=>	16918,
		60271	=>	16921,
		60272	=>	16924,
		60273	=>	16926,
		60274	=>	16929,
		60275	=>	16932,
		60276	=>	16935,
		60277	=>	16937,
		60278	=>	16940,
		60279	=>	16943,
		60280	=>	16946,
		60281	=>	16948,
		60282	=>	16951,
		60283	=>	16954,
		60284	=>	16957,
		60285	=>	16959,
		60286	=>	16962,
		60287	=>	16965,
		60288	=>	16968,
		60289	=>	16970,
		60290	=>	16973,
		60291	=>	16976,
		60292	=>	16979,
		60293	=>	16981,
		60294	=>	16984,
		60295	=>	16987,
		60296	=>	16990,
		60297	=>	16992,
		60298	=>	16995,
		60299	=>	16998,
		60300	=>	17001,
		60301	=>	17003,
		60302	=>	17006,
		60303	=>	17009,
		60304	=>	17012,
		60305	=>	17014,
		60306	=>	17017,
		60307	=>	17020,
		60308	=>	17023,
		60309	=>	17025,
		60310	=>	17028,
		60311	=>	17031,
		60312	=>	17034,
		60313	=>	17036,
		60314	=>	17039,
		60315	=>	17042,
		60316	=>	17045,
		60317	=>	17047,
		60318	=>	17050,
		60319	=>	17053,
		60320	=>	17056,
		60321	=>	17058,
		60322	=>	17061,
		60323	=>	17064,
		60324	=>	17067,
		60325	=>	17069,
		60326	=>	17072,
		60327	=>	17075,
		60328	=>	17078,
		60329	=>	17081,
		60330	=>	17083,
		60331	=>	17086,
		60332	=>	17089,
		60333	=>	17092,
		60334	=>	17094,
		60335	=>	17097,
		60336	=>	17100,
		60337	=>	17103,
		60338	=>	17105,
		60339	=>	17108,
		60340	=>	17111,
		60341	=>	17114,
		60342	=>	17116,
		60343	=>	17119,
		60344	=>	17122,
		60345	=>	17125,
		60346	=>	17127,
		60347	=>	17130,
		60348	=>	17133,
		60349	=>	17136,
		60350	=>	17138,
		60351	=>	17141,
		60352	=>	17144,
		60353	=>	17147,
		60354	=>	17150,
		60355	=>	17152,
		60356	=>	17155,
		60357	=>	17158,
		60358	=>	17161,
		60359	=>	17163,
		60360	=>	17166,
		60361	=>	17169,
		60362	=>	17172,
		60363	=>	17174,
		60364	=>	17177,
		60365	=>	17180,
		60366	=>	17183,
		60367	=>	17185,
		60368	=>	17188,
		60369	=>	17191,
		60370	=>	17194,
		60371	=>	17196,
		60372	=>	17199,
		60373	=>	17202,
		60374	=>	17205,
		60375	=>	17208,
		60376	=>	17210,
		60377	=>	17213,
		60378	=>	17216,
		60379	=>	17219,
		60380	=>	17221,
		60381	=>	17224,
		60382	=>	17227,
		60383	=>	17230,
		60384	=>	17232,
		60385	=>	17235,
		60386	=>	17238,
		60387	=>	17241,
		60388	=>	17243,
		60389	=>	17246,
		60390	=>	17249,
		60391	=>	17252,
		60392	=>	17255,
		60393	=>	17257,
		60394	=>	17260,
		60395	=>	17263,
		60396	=>	17266,
		60397	=>	17268,
		60398	=>	17271,
		60399	=>	17274,
		60400	=>	17277,
		60401	=>	17279,
		60402	=>	17282,
		60403	=>	17285,
		60404	=>	17288,
		60405	=>	17291,
		60406	=>	17293,
		60407	=>	17296,
		60408	=>	17299,
		60409	=>	17302,
		60410	=>	17304,
		60411	=>	17307,
		60412	=>	17310,
		60413	=>	17313,
		60414	=>	17315,
		60415	=>	17318,
		60416	=>	17321,
		60417	=>	17324,
		60418	=>	17327,
		60419	=>	17329,
		60420	=>	17332,
		60421	=>	17335,
		60422	=>	17338,
		60423	=>	17340,
		60424	=>	17343,
		60425	=>	17346,
		60426	=>	17349,
		60427	=>	17351,
		60428	=>	17354,
		60429	=>	17357,
		60430	=>	17360,
		60431	=>	17363,
		60432	=>	17365,
		60433	=>	17368,
		60434	=>	17371,
		60435	=>	17374,
		60436	=>	17376,
		60437	=>	17379,
		60438	=>	17382,
		60439	=>	17385,
		60440	=>	17388,
		60441	=>	17390,
		60442	=>	17393,
		60443	=>	17396,
		60444	=>	17399,
		60445	=>	17401,
		60446	=>	17404,
		60447	=>	17407,
		60448	=>	17410,
		60449	=>	17413,
		60450	=>	17415,
		60451	=>	17418,
		60452	=>	17421,
		60453	=>	17424,
		60454	=>	17426,
		60455	=>	17429,
		60456	=>	17432,
		60457	=>	17435,
		60458	=>	17437,
		60459	=>	17440,
		60460	=>	17443,
		60461	=>	17446,
		60462	=>	17449,
		60463	=>	17451,
		60464	=>	17454,
		60465	=>	17457,
		60466	=>	17460,
		60467	=>	17462,
		60468	=>	17465,
		60469	=>	17468,
		60470	=>	17471,
		60471	=>	17474,
		60472	=>	17476,
		60473	=>	17479,
		60474	=>	17482,
		60475	=>	17485,
		60476	=>	17487,
		60477	=>	17490,
		60478	=>	17493,
		60479	=>	17496,
		60480	=>	17499,
		60481	=>	17501,
		60482	=>	17504,
		60483	=>	17507,
		60484	=>	17510,
		60485	=>	17513,
		60486	=>	17515,
		60487	=>	17518,
		60488	=>	17521,
		60489	=>	17524,
		60490	=>	17526,
		60491	=>	17529,
		60492	=>	17532,
		60493	=>	17535,
		60494	=>	17538,
		60495	=>	17540,
		60496	=>	17543,
		60497	=>	17546,
		60498	=>	17549,
		60499	=>	17551,
		60500	=>	17554,
		60501	=>	17557,
		60502	=>	17560,
		60503	=>	17563,
		60504	=>	17565,
		60505	=>	17568,
		60506	=>	17571,
		60507	=>	17574,
		60508	=>	17576,
		60509	=>	17579,
		60510	=>	17582,
		60511	=>	17585,
		60512	=>	17588,
		60513	=>	17590,
		60514	=>	17593,
		60515	=>	17596,
		60516	=>	17599,
		60517	=>	17602,
		60518	=>	17604,
		60519	=>	17607,
		60520	=>	17610,
		60521	=>	17613,
		60522	=>	17615,
		60523	=>	17618,
		60524	=>	17621,
		60525	=>	17624,
		60526	=>	17627,
		60527	=>	17629,
		60528	=>	17632,
		60529	=>	17635,
		60530	=>	17638,
		60531	=>	17641,
		60532	=>	17643,
		60533	=>	17646,
		60534	=>	17649,
		60535	=>	17652,
		60536	=>	17654,
		60537	=>	17657,
		60538	=>	17660,
		60539	=>	17663,
		60540	=>	17666,
		60541	=>	17668,
		60542	=>	17671,
		60543	=>	17674,
		60544	=>	17677,
		60545	=>	17680,
		60546	=>	17682,
		60547	=>	17685,
		60548	=>	17688,
		60549	=>	17691,
		60550	=>	17694,
		60551	=>	17696,
		60552	=>	17699,
		60553	=>	17702,
		60554	=>	17705,
		60555	=>	17707,
		60556	=>	17710,
		60557	=>	17713,
		60558	=>	17716,
		60559	=>	17719,
		60560	=>	17721,
		60561	=>	17724,
		60562	=>	17727,
		60563	=>	17730,
		60564	=>	17733,
		60565	=>	17735,
		60566	=>	17738,
		60567	=>	17741,
		60568	=>	17744,
		60569	=>	17747,
		60570	=>	17749,
		60571	=>	17752,
		60572	=>	17755,
		60573	=>	17758,
		60574	=>	17761,
		60575	=>	17763,
		60576	=>	17766,
		60577	=>	17769,
		60578	=>	17772,
		60579	=>	17774,
		60580	=>	17777,
		60581	=>	17780,
		60582	=>	17783,
		60583	=>	17786,
		60584	=>	17788,
		60585	=>	17791,
		60586	=>	17794,
		60587	=>	17797,
		60588	=>	17800,
		60589	=>	17802,
		60590	=>	17805,
		60591	=>	17808,
		60592	=>	17811,
		60593	=>	17814,
		60594	=>	17816,
		60595	=>	17819,
		60596	=>	17822,
		60597	=>	17825,
		60598	=>	17828,
		60599	=>	17830,
		60600	=>	17833,
		60601	=>	17836,
		60602	=>	17839,
		60603	=>	17842,
		60604	=>	17844,
		60605	=>	17847,
		60606	=>	17850,
		60607	=>	17853,
		60608	=>	17856,
		60609	=>	17858,
		60610	=>	17861,
		60611	=>	17864,
		60612	=>	17867,
		60613	=>	17870,
		60614	=>	17872,
		60615	=>	17875,
		60616	=>	17878,
		60617	=>	17881,
		60618	=>	17884,
		60619	=>	17886,
		60620	=>	17889,
		60621	=>	17892,
		60622	=>	17895,
		60623	=>	17898,
		60624	=>	17900,
		60625	=>	17903,
		60626	=>	17906,
		60627	=>	17909,
		60628	=>	17912,
		60629	=>	17914,
		60630	=>	17917,
		60631	=>	17920,
		60632	=>	17923,
		60633	=>	17926,
		60634	=>	17928,
		60635	=>	17931,
		60636	=>	17934,
		60637	=>	17937,
		60638	=>	17940,
		60639	=>	17942,
		60640	=>	17945,
		60641	=>	17948,
		60642	=>	17951,
		60643	=>	17954,
		60644	=>	17956,
		60645	=>	17959,
		60646	=>	17962,
		60647	=>	17965,
		60648	=>	17968,
		60649	=>	17970,
		60650	=>	17973,
		60651	=>	17976,
		60652	=>	17979,
		60653	=>	17982,
		60654	=>	17984,
		60655	=>	17987,
		60656	=>	17990,
		60657	=>	17993,
		60658	=>	17996,
		60659	=>	17998,
		60660	=>	18001,
		60661	=>	18004,
		60662	=>	18007,
		60663	=>	18010,
		60664	=>	18012,
		60665	=>	18015,
		60666	=>	18018,
		60667	=>	18021,
		60668	=>	18024,
		60669	=>	18026,
		60670	=>	18029,
		60671	=>	18032,
		60672	=>	18035,
		60673	=>	18038,
		60674	=>	18040,
		60675	=>	18043,
		60676	=>	18046,
		60677	=>	18049,
		60678	=>	18052,
		60679	=>	18055,
		60680	=>	18057,
		60681	=>	18060,
		60682	=>	18063,
		60683	=>	18066,
		60684	=>	18069,
		60685	=>	18071,
		60686	=>	18074,
		60687	=>	18077,
		60688	=>	18080,
		60689	=>	18083,
		60690	=>	18085,
		60691	=>	18088,
		60692	=>	18091,
		60693	=>	18094,
		60694	=>	18097,
		60695	=>	18099,
		60696	=>	18102,
		60697	=>	18105,
		60698	=>	18108,
		60699	=>	18111,
		60700	=>	18113,
		60701	=>	18116,
		60702	=>	18119,
		60703	=>	18122,
		60704	=>	18125,
		60705	=>	18128,
		60706	=>	18130,
		60707	=>	18133,
		60708	=>	18136,
		60709	=>	18139,
		60710	=>	18142,
		60711	=>	18144,
		60712	=>	18147,
		60713	=>	18150,
		60714	=>	18153,
		60715	=>	18156,
		60716	=>	18158,
		60717	=>	18161,
		60718	=>	18164,
		60719	=>	18167,
		60720	=>	18170,
		60721	=>	18173,
		60722	=>	18175,
		60723	=>	18178,
		60724	=>	18181,
		60725	=>	18184,
		60726	=>	18187,
		60727	=>	18189,
		60728	=>	18192,
		60729	=>	18195,
		60730	=>	18198,
		60731	=>	18201,
		60732	=>	18203,
		60733	=>	18206,
		60734	=>	18209,
		60735	=>	18212,
		60736	=>	18215,
		60737	=>	18218,
		60738	=>	18220,
		60739	=>	18223,
		60740	=>	18226,
		60741	=>	18229,
		60742	=>	18232,
		60743	=>	18234,
		60744	=>	18237,
		60745	=>	18240,
		60746	=>	18243,
		60747	=>	18246,
		60748	=>	18249,
		60749	=>	18251,
		60750	=>	18254,
		60751	=>	18257,
		60752	=>	18260,
		60753	=>	18263,
		60754	=>	18265,
		60755	=>	18268,
		60756	=>	18271,
		60757	=>	18274,
		60758	=>	18277,
		60759	=>	18280,
		60760	=>	18282,
		60761	=>	18285,
		60762	=>	18288,
		60763	=>	18291,
		60764	=>	18294,
		60765	=>	18296,
		60766	=>	18299,
		60767	=>	18302,
		60768	=>	18305,
		60769	=>	18308,
		60770	=>	18311,
		60771	=>	18313,
		60772	=>	18316,
		60773	=>	18319,
		60774	=>	18322,
		60775	=>	18325,
		60776	=>	18327,
		60777	=>	18330,
		60778	=>	18333,
		60779	=>	18336,
		60780	=>	18339,
		60781	=>	18342,
		60782	=>	18344,
		60783	=>	18347,
		60784	=>	18350,
		60785	=>	18353,
		60786	=>	18356,
		60787	=>	18358,
		60788	=>	18361,
		60789	=>	18364,
		60790	=>	18367,
		60791	=>	18370,
		60792	=>	18373,
		60793	=>	18375,
		60794	=>	18378,
		60795	=>	18381,
		60796	=>	18384,
		60797	=>	18387,
		60798	=>	18389,
		60799	=>	18392,
		60800	=>	18395,
		60801	=>	18398,
		60802	=>	18401,
		60803	=>	18404,
		60804	=>	18406,
		60805	=>	18409,
		60806	=>	18412,
		60807	=>	18415,
		60808	=>	18418,
		60809	=>	18421,
		60810	=>	18423,
		60811	=>	18426,
		60812	=>	18429,
		60813	=>	18432,
		60814	=>	18435,
		60815	=>	18438,
		60816	=>	18440,
		60817	=>	18443,
		60818	=>	18446,
		60819	=>	18449,
		60820	=>	18452,
		60821	=>	18454,
		60822	=>	18457,
		60823	=>	18460,
		60824	=>	18463,
		60825	=>	18466,
		60826	=>	18469,
		60827	=>	18471,
		60828	=>	18474,
		60829	=>	18477,
		60830	=>	18480,
		60831	=>	18483,
		60832	=>	18486,
		60833	=>	18488,
		60834	=>	18491,
		60835	=>	18494,
		60836	=>	18497,
		60837	=>	18500,
		60838	=>	18503,
		60839	=>	18505,
		60840	=>	18508,
		60841	=>	18511,
		60842	=>	18514,
		60843	=>	18517,
		60844	=>	18519,
		60845	=>	18522,
		60846	=>	18525,
		60847	=>	18528,
		60848	=>	18531,
		60849	=>	18534,
		60850	=>	18536,
		60851	=>	18539,
		60852	=>	18542,
		60853	=>	18545,
		60854	=>	18548,
		60855	=>	18551,
		60856	=>	18553,
		60857	=>	18556,
		60858	=>	18559,
		60859	=>	18562,
		60860	=>	18565,
		60861	=>	18568,
		60862	=>	18570,
		60863	=>	18573,
		60864	=>	18576,
		60865	=>	18579,
		60866	=>	18582,
		60867	=>	18585,
		60868	=>	18587,
		60869	=>	18590,
		60870	=>	18593,
		60871	=>	18596,
		60872	=>	18599,
		60873	=>	18602,
		60874	=>	18604,
		60875	=>	18607,
		60876	=>	18610,
		60877	=>	18613,
		60878	=>	18616,
		60879	=>	18619,
		60880	=>	18621,
		60881	=>	18624,
		60882	=>	18627,
		60883	=>	18630,
		60884	=>	18633,
		60885	=>	18636,
		60886	=>	18638,
		60887	=>	18641,
		60888	=>	18644,
		60889	=>	18647,
		60890	=>	18650,
		60891	=>	18653,
		60892	=>	18655,
		60893	=>	18658,
		60894	=>	18661,
		60895	=>	18664,
		60896	=>	18667,
		60897	=>	18670,
		60898	=>	18672,
		60899	=>	18675,
		60900	=>	18678,
		60901	=>	18681,
		60902	=>	18684,
		60903	=>	18687,
		60904	=>	18689,
		60905	=>	18692,
		60906	=>	18695,
		60907	=>	18698,
		60908	=>	18701,
		60909	=>	18704,
		60910	=>	18706,
		60911	=>	18709,
		60912	=>	18712,
		60913	=>	18715,
		60914	=>	18718,
		60915	=>	18721,
		60916	=>	18724,
		60917	=>	18726,
		60918	=>	18729,
		60919	=>	18732,
		60920	=>	18735,
		60921	=>	18738,
		60922	=>	18741,
		60923	=>	18743,
		60924	=>	18746,
		60925	=>	18749,
		60926	=>	18752,
		60927	=>	18755,
		60928	=>	18758,
		60929	=>	18760,
		60930	=>	18763,
		60931	=>	18766,
		60932	=>	18769,
		60933	=>	18772,
		60934	=>	18775,
		60935	=>	18777,
		60936	=>	18780,
		60937	=>	18783,
		60938	=>	18786,
		60939	=>	18789,
		60940	=>	18792,
		60941	=>	18795,
		60942	=>	18797,
		60943	=>	18800,
		60944	=>	18803,
		60945	=>	18806,
		60946	=>	18809,
		60947	=>	18812,
		60948	=>	18814,
		60949	=>	18817,
		60950	=>	18820,
		60951	=>	18823,
		60952	=>	18826,
		60953	=>	18829,
		60954	=>	18831,
		60955	=>	18834,
		60956	=>	18837,
		60957	=>	18840,
		60958	=>	18843,
		60959	=>	18846,
		60960	=>	18849,
		60961	=>	18851,
		60962	=>	18854,
		60963	=>	18857,
		60964	=>	18860,
		60965	=>	18863,
		60966	=>	18866,
		60967	=>	18868,
		60968	=>	18871,
		60969	=>	18874,
		60970	=>	18877,
		60971	=>	18880,
		60972	=>	18883,
		60973	=>	18886,
		60974	=>	18888,
		60975	=>	18891,
		60976	=>	18894,
		60977	=>	18897,
		60978	=>	18900,
		60979	=>	18903,
		60980	=>	18905,
		60981	=>	18908,
		60982	=>	18911,
		60983	=>	18914,
		60984	=>	18917,
		60985	=>	18920,
		60986	=>	18923,
		60987	=>	18925,
		60988	=>	18928,
		60989	=>	18931,
		60990	=>	18934,
		60991	=>	18937,
		60992	=>	18940,
		60993	=>	18942,
		60994	=>	18945,
		60995	=>	18948,
		60996	=>	18951,
		60997	=>	18954,
		60998	=>	18957,
		60999	=>	18960,
		61000	=>	18962,
		61001	=>	18965,
		61002	=>	18968,
		61003	=>	18971,
		61004	=>	18974,
		61005	=>	18977,
		61006	=>	18979,
		61007	=>	18982,
		61008	=>	18985,
		61009	=>	18988,
		61010	=>	18991,
		61011	=>	18994,
		61012	=>	18997,
		61013	=>	18999,
		61014	=>	19002,
		61015	=>	19005,
		61016	=>	19008,
		61017	=>	19011,
		61018	=>	19014,
		61019	=>	19017,
		61020	=>	19019,
		61021	=>	19022,
		61022	=>	19025,
		61023	=>	19028,
		61024	=>	19031,
		61025	=>	19034,
		61026	=>	19037,
		61027	=>	19039,
		61028	=>	19042,
		61029	=>	19045,
		61030	=>	19048,
		61031	=>	19051,
		61032	=>	19054,
		61033	=>	19056,
		61034	=>	19059,
		61035	=>	19062,
		61036	=>	19065,
		61037	=>	19068,
		61038	=>	19071,
		61039	=>	19074,
		61040	=>	19076,
		61041	=>	19079,
		61042	=>	19082,
		61043	=>	19085,
		61044	=>	19088,
		61045	=>	19091,
		61046	=>	19094,
		61047	=>	19096,
		61048	=>	19099,
		61049	=>	19102,
		61050	=>	19105,
		61051	=>	19108,
		61052	=>	19111,
		61053	=>	19114,
		61054	=>	19116,
		61055	=>	19119,
		61056	=>	19122,
		61057	=>	19125,
		61058	=>	19128,
		61059	=>	19131,
		61060	=>	19134,
		61061	=>	19136,
		61062	=>	19139,
		61063	=>	19142,
		61064	=>	19145,
		61065	=>	19148,
		61066	=>	19151,
		61067	=>	19154,
		61068	=>	19156,
		61069	=>	19159,
		61070	=>	19162,
		61071	=>	19165,
		61072	=>	19168,
		61073	=>	19171,
		61074	=>	19174,
		61075	=>	19176,
		61076	=>	19179,
		61077	=>	19182,
		61078	=>	19185,
		61079	=>	19188,
		61080	=>	19191,
		61081	=>	19194,
		61082	=>	19196,
		61083	=>	19199,
		61084	=>	19202,
		61085	=>	19205,
		61086	=>	19208,
		61087	=>	19211,
		61088	=>	19214,
		61089	=>	19216,
		61090	=>	19219,
		61091	=>	19222,
		61092	=>	19225,
		61093	=>	19228,
		61094	=>	19231,
		61095	=>	19234,
		61096	=>	19236,
		61097	=>	19239,
		61098	=>	19242,
		61099	=>	19245,
		61100	=>	19248,
		61101	=>	19251,
		61102	=>	19254,
		61103	=>	19257,
		61104	=>	19259,
		61105	=>	19262,
		61106	=>	19265,
		61107	=>	19268,
		61108	=>	19271,
		61109	=>	19274,
		61110	=>	19277,
		61111	=>	19279,
		61112	=>	19282,
		61113	=>	19285,
		61114	=>	19288,
		61115	=>	19291,
		61116	=>	19294,
		61117	=>	19297,
		61118	=>	19299,
		61119	=>	19302,
		61120	=>	19305,
		61121	=>	19308,
		61122	=>	19311,
		61123	=>	19314,
		61124	=>	19317,
		61125	=>	19320,
		61126	=>	19322,
		61127	=>	19325,
		61128	=>	19328,
		61129	=>	19331,
		61130	=>	19334,
		61131	=>	19337,
		61132	=>	19340,
		61133	=>	19342,
		61134	=>	19345,
		61135	=>	19348,
		61136	=>	19351,
		61137	=>	19354,
		61138	=>	19357,
		61139	=>	19360,
		61140	=>	19363,
		61141	=>	19365,
		61142	=>	19368,
		61143	=>	19371,
		61144	=>	19374,
		61145	=>	19377,
		61146	=>	19380,
		61147	=>	19383,
		61148	=>	19385,
		61149	=>	19388,
		61150	=>	19391,
		61151	=>	19394,
		61152	=>	19397,
		61153	=>	19400,
		61154	=>	19403,
		61155	=>	19406,
		61156	=>	19408,
		61157	=>	19411,
		61158	=>	19414,
		61159	=>	19417,
		61160	=>	19420,
		61161	=>	19423,
		61162	=>	19426,
		61163	=>	19428,
		61164	=>	19431,
		61165	=>	19434,
		61166	=>	19437,
		61167	=>	19440,
		61168	=>	19443,
		61169	=>	19446,
		61170	=>	19449,
		61171	=>	19451,
		61172	=>	19454,
		61173	=>	19457,
		61174	=>	19460,
		61175	=>	19463,
		61176	=>	19466,
		61177	=>	19469,
		61178	=>	19472,
		61179	=>	19474,
		61180	=>	19477,
		61181	=>	19480,
		61182	=>	19483,
		61183	=>	19486,
		61184	=>	19489,
		61185	=>	19492,
		61186	=>	19494,
		61187	=>	19497,
		61188	=>	19500,
		61189	=>	19503,
		61190	=>	19506,
		61191	=>	19509,
		61192	=>	19512,
		61193	=>	19515,
		61194	=>	19517,
		61195	=>	19520,
		61196	=>	19523,
		61197	=>	19526,
		61198	=>	19529,
		61199	=>	19532,
		61200	=>	19535,
		61201	=>	19538,
		61202	=>	19540,
		61203	=>	19543,
		61204	=>	19546,
		61205	=>	19549,
		61206	=>	19552,
		61207	=>	19555,
		61208	=>	19558,
		61209	=>	19561,
		61210	=>	19563,
		61211	=>	19566,
		61212	=>	19569,
		61213	=>	19572,
		61214	=>	19575,
		61215	=>	19578,
		61216	=>	19581,
		61217	=>	19584,
		61218	=>	19586,
		61219	=>	19589,
		61220	=>	19592,
		61221	=>	19595,
		61222	=>	19598,
		61223	=>	19601,
		61224	=>	19604,
		61225	=>	19607,
		61226	=>	19609,
		61227	=>	19612,
		61228	=>	19615,
		61229	=>	19618,
		61230	=>	19621,
		61231	=>	19624,
		61232	=>	19627,
		61233	=>	19630,
		61234	=>	19633,
		61235	=>	19635,
		61236	=>	19638,
		61237	=>	19641,
		61238	=>	19644,
		61239	=>	19647,
		61240	=>	19650,
		61241	=>	19653,
		61242	=>	19656,
		61243	=>	19658,
		61244	=>	19661,
		61245	=>	19664,
		61246	=>	19667,
		61247	=>	19670,
		61248	=>	19673,
		61249	=>	19676,
		61250	=>	19679,
		61251	=>	19681,
		61252	=>	19684,
		61253	=>	19687,
		61254	=>	19690,
		61255	=>	19693,
		61256	=>	19696,
		61257	=>	19699,
		61258	=>	19702,
		61259	=>	19704,
		61260	=>	19707,
		61261	=>	19710,
		61262	=>	19713,
		61263	=>	19716,
		61264	=>	19719,
		61265	=>	19722,
		61266	=>	19725,
		61267	=>	19728,
		61268	=>	19730,
		61269	=>	19733,
		61270	=>	19736,
		61271	=>	19739,
		61272	=>	19742,
		61273	=>	19745,
		61274	=>	19748,
		61275	=>	19751,
		61276	=>	19753,
		61277	=>	19756,
		61278	=>	19759,
		61279	=>	19762,
		61280	=>	19765,
		61281	=>	19768,
		61282	=>	19771,
		61283	=>	19774,
		61284	=>	19777,
		61285	=>	19779,
		61286	=>	19782,
		61287	=>	19785,
		61288	=>	19788,
		61289	=>	19791,
		61290	=>	19794,
		61291	=>	19797,
		61292	=>	19800,
		61293	=>	19803,
		61294	=>	19805,
		61295	=>	19808,
		61296	=>	19811,
		61297	=>	19814,
		61298	=>	19817,
		61299	=>	19820,
		61300	=>	19823,
		61301	=>	19826,
		61302	=>	19828,
		61303	=>	19831,
		61304	=>	19834,
		61305	=>	19837,
		61306	=>	19840,
		61307	=>	19843,
		61308	=>	19846,
		61309	=>	19849,
		61310	=>	19852,
		61311	=>	19854,
		61312	=>	19857,
		61313	=>	19860,
		61314	=>	19863,
		61315	=>	19866,
		61316	=>	19869,
		61317	=>	19872,
		61318	=>	19875,
		61319	=>	19878,
		61320	=>	19880,
		61321	=>	19883,
		61322	=>	19886,
		61323	=>	19889,
		61324	=>	19892,
		61325	=>	19895,
		61326	=>	19898,
		61327	=>	19901,
		61328	=>	19904,
		61329	=>	19906,
		61330	=>	19909,
		61331	=>	19912,
		61332	=>	19915,
		61333	=>	19918,
		61334	=>	19921,
		61335	=>	19924,
		61336	=>	19927,
		61337	=>	19930,
		61338	=>	19932,
		61339	=>	19935,
		61340	=>	19938,
		61341	=>	19941,
		61342	=>	19944,
		61343	=>	19947,
		61344	=>	19950,
		61345	=>	19953,
		61346	=>	19956,
		61347	=>	19958,
		61348	=>	19961,
		61349	=>	19964,
		61350	=>	19967,
		61351	=>	19970,
		61352	=>	19973,
		61353	=>	19976,
		61354	=>	19979,
		61355	=>	19982,
		61356	=>	19985,
		61357	=>	19987,
		61358	=>	19990,
		61359	=>	19993,
		61360	=>	19996,
		61361	=>	19999,
		61362	=>	20002,
		61363	=>	20005,
		61364	=>	20008,
		61365	=>	20011,
		61366	=>	20013,
		61367	=>	20016,
		61368	=>	20019,
		61369	=>	20022,
		61370	=>	20025,
		61371	=>	20028,
		61372	=>	20031,
		61373	=>	20034,
		61374	=>	20037,
		61375	=>	20040,
		61376	=>	20042,
		61377	=>	20045,
		61378	=>	20048,
		61379	=>	20051,
		61380	=>	20054,
		61381	=>	20057,
		61382	=>	20060,
		61383	=>	20063,
		61384	=>	20066,
		61385	=>	20068,
		61386	=>	20071,
		61387	=>	20074,
		61388	=>	20077,
		61389	=>	20080,
		61390	=>	20083,
		61391	=>	20086,
		61392	=>	20089,
		61393	=>	20092,
		61394	=>	20095,
		61395	=>	20097,
		61396	=>	20100,
		61397	=>	20103,
		61398	=>	20106,
		61399	=>	20109,
		61400	=>	20112,
		61401	=>	20115,
		61402	=>	20118,
		61403	=>	20121,
		61404	=>	20124,
		61405	=>	20126,
		61406	=>	20129,
		61407	=>	20132,
		61408	=>	20135,
		61409	=>	20138,
		61410	=>	20141,
		61411	=>	20144,
		61412	=>	20147,
		61413	=>	20150,
		61414	=>	20152,
		61415	=>	20155,
		61416	=>	20158,
		61417	=>	20161,
		61418	=>	20164,
		61419	=>	20167,
		61420	=>	20170,
		61421	=>	20173,
		61422	=>	20176,
		61423	=>	20179,
		61424	=>	20181,
		61425	=>	20184,
		61426	=>	20187,
		61427	=>	20190,
		61428	=>	20193,
		61429	=>	20196,
		61430	=>	20199,
		61431	=>	20202,
		61432	=>	20205,
		61433	=>	20208,
		61434	=>	20211,
		61435	=>	20213,
		61436	=>	20216,
		61437	=>	20219,
		61438	=>	20222,
		61439	=>	20225,
		61440	=>	20228,
		61441	=>	20231,
		61442	=>	20234,
		61443	=>	20237,
		61444	=>	20240,
		61445	=>	20242,
		61446	=>	20245,
		61447	=>	20248,
		61448	=>	20251,
		61449	=>	20254,
		61450	=>	20257,
		61451	=>	20260,
		61452	=>	20263,
		61453	=>	20266,
		61454	=>	20269,
		61455	=>	20271,
		61456	=>	20274,
		61457	=>	20277,
		61458	=>	20280,
		61459	=>	20283,
		61460	=>	20286,
		61461	=>	20289,
		61462	=>	20292,
		61463	=>	20295,
		61464	=>	20298,
		61465	=>	20301,
		61466	=>	20303,
		61467	=>	20306,
		61468	=>	20309,
		61469	=>	20312,
		61470	=>	20315,
		61471	=>	20318,
		61472	=>	20321,
		61473	=>	20324,
		61474	=>	20327,
		61475	=>	20330,
		61476	=>	20332,
		61477	=>	20335,
		61478	=>	20338,
		61479	=>	20341,
		61480	=>	20344,
		61481	=>	20347,
		61482	=>	20350,
		61483	=>	20353,
		61484	=>	20356,
		61485	=>	20359,
		61486	=>	20362,
		61487	=>	20364,
		61488	=>	20367,
		61489	=>	20370,
		61490	=>	20373,
		61491	=>	20376,
		61492	=>	20379,
		61493	=>	20382,
		61494	=>	20385,
		61495	=>	20388,
		61496	=>	20391,
		61497	=>	20394,
		61498	=>	20396,
		61499	=>	20399,
		61500	=>	20402,
		61501	=>	20405,
		61502	=>	20408,
		61503	=>	20411,
		61504	=>	20414,
		61505	=>	20417,
		61506	=>	20420,
		61507	=>	20423,
		61508	=>	20426,
		61509	=>	20428,
		61510	=>	20431,
		61511	=>	20434,
		61512	=>	20437,
		61513	=>	20440,
		61514	=>	20443,
		61515	=>	20446,
		61516	=>	20449,
		61517	=>	20452,
		61518	=>	20455,
		61519	=>	20458,
		61520	=>	20460,
		61521	=>	20463,
		61522	=>	20466,
		61523	=>	20469,
		61524	=>	20472,
		61525	=>	20475,
		61526	=>	20478,
		61527	=>	20481,
		61528	=>	20484,
		61529	=>	20487,
		61530	=>	20490,
		61531	=>	20493,
		61532	=>	20495,
		61533	=>	20498,
		61534	=>	20501,
		61535	=>	20504,
		61536	=>	20507,
		61537	=>	20510,
		61538	=>	20513,
		61539	=>	20516,
		61540	=>	20519,
		61541	=>	20522,
		61542	=>	20525,
		61543	=>	20527,
		61544	=>	20530,
		61545	=>	20533,
		61546	=>	20536,
		61547	=>	20539,
		61548	=>	20542,
		61549	=>	20545,
		61550	=>	20548,
		61551	=>	20551,
		61552	=>	20554,
		61553	=>	20557,
		61554	=>	20560,
		61555	=>	20562,
		61556	=>	20565,
		61557	=>	20568,
		61558	=>	20571,
		61559	=>	20574,
		61560	=>	20577,
		61561	=>	20580,
		61562	=>	20583,
		61563	=>	20586,
		61564	=>	20589,
		61565	=>	20592,
		61566	=>	20595,
		61567	=>	20597,
		61568	=>	20600,
		61569	=>	20603,
		61570	=>	20606,
		61571	=>	20609,
		61572	=>	20612,
		61573	=>	20615,
		61574	=>	20618,
		61575	=>	20621,
		61576	=>	20624,
		61577	=>	20627,
		61578	=>	20630,
		61579	=>	20632,
		61580	=>	20635,
		61581	=>	20638,
		61582	=>	20641,
		61583	=>	20644,
		61584	=>	20647,
		61585	=>	20650,
		61586	=>	20653,
		61587	=>	20656,
		61588	=>	20659,
		61589	=>	20662,
		61590	=>	20665,
		61591	=>	20667,
		61592	=>	20670,
		61593	=>	20673,
		61594	=>	20676,
		61595	=>	20679,
		61596	=>	20682,
		61597	=>	20685,
		61598	=>	20688,
		61599	=>	20691,
		61600	=>	20694,
		61601	=>	20697,
		61602	=>	20700,
		61603	=>	20703,
		61604	=>	20705,
		61605	=>	20708,
		61606	=>	20711,
		61607	=>	20714,
		61608	=>	20717,
		61609	=>	20720,
		61610	=>	20723,
		61611	=>	20726,
		61612	=>	20729,
		61613	=>	20732,
		61614	=>	20735,
		61615	=>	20738,
		61616	=>	20741,
		61617	=>	20743,
		61618	=>	20746,
		61619	=>	20749,
		61620	=>	20752,
		61621	=>	20755,
		61622	=>	20758,
		61623	=>	20761,
		61624	=>	20764,
		61625	=>	20767,
		61626	=>	20770,
		61627	=>	20773,
		61628	=>	20776,
		61629	=>	20779,
		61630	=>	20781,
		61631	=>	20784,
		61632	=>	20787,
		61633	=>	20790,
		61634	=>	20793,
		61635	=>	20796,
		61636	=>	20799,
		61637	=>	20802,
		61638	=>	20805,
		61639	=>	20808,
		61640	=>	20811,
		61641	=>	20814,
		61642	=>	20817,
		61643	=>	20819,
		61644	=>	20822,
		61645	=>	20825,
		61646	=>	20828,
		61647	=>	20831,
		61648	=>	20834,
		61649	=>	20837,
		61650	=>	20840,
		61651	=>	20843,
		61652	=>	20846,
		61653	=>	20849,
		61654	=>	20852,
		61655	=>	20855,
		61656	=>	20857,
		61657	=>	20860,
		61658	=>	20863,
		61659	=>	20866,
		61660	=>	20869,
		61661	=>	20872,
		61662	=>	20875,
		61663	=>	20878,
		61664	=>	20881,
		61665	=>	20884,
		61666	=>	20887,
		61667	=>	20890,
		61668	=>	20893,
		61669	=>	20896,
		61670	=>	20898,
		61671	=>	20901,
		61672	=>	20904,
		61673	=>	20907,
		61674	=>	20910,
		61675	=>	20913,
		61676	=>	20916,
		61677	=>	20919,
		61678	=>	20922,
		61679	=>	20925,
		61680	=>	20928,
		61681	=>	20931,
		61682	=>	20934,
		61683	=>	20937,
		61684	=>	20939,
		61685	=>	20942,
		61686	=>	20945,
		61687	=>	20948,
		61688	=>	20951,
		61689	=>	20954,
		61690	=>	20957,
		61691	=>	20960,
		61692	=>	20963,
		61693	=>	20966,
		61694	=>	20969,
		61695	=>	20972,
		61696	=>	20975,
		61697	=>	20978,
		61698	=>	20981,
		61699	=>	20983,
		61700	=>	20986,
		61701	=>	20989,
		61702	=>	20992,
		61703	=>	20995,
		61704	=>	20998,
		61705	=>	21001,
		61706	=>	21004,
		61707	=>	21007,
		61708	=>	21010,
		61709	=>	21013,
		61710	=>	21016,
		61711	=>	21019,
		61712	=>	21022,
		61713	=>	21024,
		61714	=>	21027,
		61715	=>	21030,
		61716	=>	21033,
		61717	=>	21036,
		61718	=>	21039,
		61719	=>	21042,
		61720	=>	21045,
		61721	=>	21048,
		61722	=>	21051,
		61723	=>	21054,
		61724	=>	21057,
		61725	=>	21060,
		61726	=>	21063,
		61727	=>	21066,
		61728	=>	21068,
		61729	=>	21071,
		61730	=>	21074,
		61731	=>	21077,
		61732	=>	21080,
		61733	=>	21083,
		61734	=>	21086,
		61735	=>	21089,
		61736	=>	21092,
		61737	=>	21095,
		61738	=>	21098,
		61739	=>	21101,
		61740	=>	21104,
		61741	=>	21107,
		61742	=>	21110,
		61743	=>	21113,
		61744	=>	21115,
		61745	=>	21118,
		61746	=>	21121,
		61747	=>	21124,
		61748	=>	21127,
		61749	=>	21130,
		61750	=>	21133,
		61751	=>	21136,
		61752	=>	21139,
		61753	=>	21142,
		61754	=>	21145,
		61755	=>	21148,
		61756	=>	21151,
		61757	=>	21154,
		61758	=>	21157,
		61759	=>	21160,
		61760	=>	21162,
		61761	=>	21165,
		61762	=>	21168,
		61763	=>	21171,
		61764	=>	21174,
		61765	=>	21177,
		61766	=>	21180,
		61767	=>	21183,
		61768	=>	21186,
		61769	=>	21189,
		61770	=>	21192,
		61771	=>	21195,
		61772	=>	21198,
		61773	=>	21201,
		61774	=>	21204,
		61775	=>	21207,
		61776	=>	21209,
		61777	=>	21212,
		61778	=>	21215,
		61779	=>	21218,
		61780	=>	21221,
		61781	=>	21224,
		61782	=>	21227,
		61783	=>	21230,
		61784	=>	21233,
		61785	=>	21236,
		61786	=>	21239,
		61787	=>	21242,
		61788	=>	21245,
		61789	=>	21248,
		61790	=>	21251,
		61791	=>	21254,
		61792	=>	21257,
		61793	=>	21259,
		61794	=>	21262,
		61795	=>	21265,
		61796	=>	21268,
		61797	=>	21271,
		61798	=>	21274,
		61799	=>	21277,
		61800	=>	21280,
		61801	=>	21283,
		61802	=>	21286,
		61803	=>	21289,
		61804	=>	21292,
		61805	=>	21295,
		61806	=>	21298,
		61807	=>	21301,
		61808	=>	21304,
		61809	=>	21307,
		61810	=>	21309,
		61811	=>	21312,
		61812	=>	21315,
		61813	=>	21318,
		61814	=>	21321,
		61815	=>	21324,
		61816	=>	21327,
		61817	=>	21330,
		61818	=>	21333,
		61819	=>	21336,
		61820	=>	21339,
		61821	=>	21342,
		61822	=>	21345,
		61823	=>	21348,
		61824	=>	21351,
		61825	=>	21354,
		61826	=>	21357,
		61827	=>	21360,
		61828	=>	21362,
		61829	=>	21365,
		61830	=>	21368,
		61831	=>	21371,
		61832	=>	21374,
		61833	=>	21377,
		61834	=>	21380,
		61835	=>	21383,
		61836	=>	21386,
		61837	=>	21389,
		61838	=>	21392,
		61839	=>	21395,
		61840	=>	21398,
		61841	=>	21401,
		61842	=>	21404,
		61843	=>	21407,
		61844	=>	21410,
		61845	=>	21413,
		61846	=>	21415,
		61847	=>	21418,
		61848	=>	21421,
		61849	=>	21424,
		61850	=>	21427,
		61851	=>	21430,
		61852	=>	21433,
		61853	=>	21436,
		61854	=>	21439,
		61855	=>	21442,
		61856	=>	21445,
		61857	=>	21448,
		61858	=>	21451,
		61859	=>	21454,
		61860	=>	21457,
		61861	=>	21460,
		61862	=>	21463,
		61863	=>	21466,
		61864	=>	21469,
		61865	=>	21472,
		61866	=>	21474,
		61867	=>	21477,
		61868	=>	21480,
		61869	=>	21483,
		61870	=>	21486,
		61871	=>	21489,
		61872	=>	21492,
		61873	=>	21495,
		61874	=>	21498,
		61875	=>	21501,
		61876	=>	21504,
		61877	=>	21507,
		61878	=>	21510,
		61879	=>	21513,
		61880	=>	21516,
		61881	=>	21519,
		61882	=>	21522,
		61883	=>	21525,
		61884	=>	21528,
		61885	=>	21531,
		61886	=>	21533,
		61887	=>	21536,
		61888	=>	21539,
		61889	=>	21542,
		61890	=>	21545,
		61891	=>	21548,
		61892	=>	21551,
		61893	=>	21554,
		61894	=>	21557,
		61895	=>	21560,
		61896	=>	21563,
		61897	=>	21566,
		61898	=>	21569,
		61899	=>	21572,
		61900	=>	21575,
		61901	=>	21578,
		61902	=>	21581,
		61903	=>	21584,
		61904	=>	21587,
		61905	=>	21590,
		61906	=>	21593,
		61907	=>	21595,
		61908	=>	21598,
		61909	=>	21601,
		61910	=>	21604,
		61911	=>	21607,
		61912	=>	21610,
		61913	=>	21613,
		61914	=>	21616,
		61915	=>	21619,
		61916	=>	21622,
		61917	=>	21625,
		61918	=>	21628,
		61919	=>	21631,
		61920	=>	21634,
		61921	=>	21637,
		61922	=>	21640,
		61923	=>	21643,
		61924	=>	21646,
		61925	=>	21649,
		61926	=>	21652,
		61927	=>	21655,
		61928	=>	21658,
		61929	=>	21660,
		61930	=>	21663,
		61931	=>	21666,
		61932	=>	21669,
		61933	=>	21672,
		61934	=>	21675,
		61935	=>	21678,
		61936	=>	21681,
		61937	=>	21684,
		61938	=>	21687,
		61939	=>	21690,
		61940	=>	21693,
		61941	=>	21696,
		61942	=>	21699,
		61943	=>	21702,
		61944	=>	21705,
		61945	=>	21708,
		61946	=>	21711,
		61947	=>	21714,
		61948	=>	21717,
		61949	=>	21720,
		61950	=>	21723,
		61951	=>	21726,
		61952	=>	21728,
		61953	=>	21731,
		61954	=>	21734,
		61955	=>	21737,
		61956	=>	21740,
		61957	=>	21743,
		61958	=>	21746,
		61959	=>	21749,
		61960	=>	21752,
		61961	=>	21755,
		61962	=>	21758,
		61963	=>	21761,
		61964	=>	21764,
		61965	=>	21767,
		61966	=>	21770,
		61967	=>	21773,
		61968	=>	21776,
		61969	=>	21779,
		61970	=>	21782,
		61971	=>	21785,
		61972	=>	21788,
		61973	=>	21791,
		61974	=>	21794,
		61975	=>	21797,
		61976	=>	21799,
		61977	=>	21802,
		61978	=>	21805,
		61979	=>	21808,
		61980	=>	21811,
		61981	=>	21814,
		61982	=>	21817,
		61983	=>	21820,
		61984	=>	21823,
		61985	=>	21826,
		61986	=>	21829,
		61987	=>	21832,
		61988	=>	21835,
		61989	=>	21838,
		61990	=>	21841,
		61991	=>	21844,
		61992	=>	21847,
		61993	=>	21850,
		61994	=>	21853,
		61995	=>	21856,
		61996	=>	21859,
		61997	=>	21862,
		61998	=>	21865,
		61999	=>	21868,
		62000	=>	21871,
		62001	=>	21874,
		62002	=>	21876,
		62003	=>	21879,
		62004	=>	21882,
		62005	=>	21885,
		62006	=>	21888,
		62007	=>	21891,
		62008	=>	21894,
		62009	=>	21897,
		62010	=>	21900,
		62011	=>	21903,
		62012	=>	21906,
		62013	=>	21909,
		62014	=>	21912,
		62015	=>	21915,
		62016	=>	21918,
		62017	=>	21921,
		62018	=>	21924,
		62019	=>	21927,
		62020	=>	21930,
		62021	=>	21933,
		62022	=>	21936,
		62023	=>	21939,
		62024	=>	21942,
		62025	=>	21945,
		62026	=>	21948,
		62027	=>	21951,
		62028	=>	21954,
		62029	=>	21957,
		62030	=>	21959,
		62031	=>	21962,
		62032	=>	21965,
		62033	=>	21968,
		62034	=>	21971,
		62035	=>	21974,
		62036	=>	21977,
		62037	=>	21980,
		62038	=>	21983,
		62039	=>	21986,
		62040	=>	21989,
		62041	=>	21992,
		62042	=>	21995,
		62043	=>	21998,
		62044	=>	22001,
		62045	=>	22004,
		62046	=>	22007,
		62047	=>	22010,
		62048	=>	22013,
		62049	=>	22016,
		62050	=>	22019,
		62051	=>	22022,
		62052	=>	22025,
		62053	=>	22028,
		62054	=>	22031,
		62055	=>	22034,
		62056	=>	22037,
		62057	=>	22040,
		62058	=>	22043,
		62059	=>	22046,
		62060	=>	22049,
		62061	=>	22051,
		62062	=>	22054,
		62063	=>	22057,
		62064	=>	22060,
		62065	=>	22063,
		62066	=>	22066,
		62067	=>	22069,
		62068	=>	22072,
		62069	=>	22075,
		62070	=>	22078,
		62071	=>	22081,
		62072	=>	22084,
		62073	=>	22087,
		62074	=>	22090,
		62075	=>	22093,
		62076	=>	22096,
		62077	=>	22099,
		62078	=>	22102,
		62079	=>	22105,
		62080	=>	22108,
		62081	=>	22111,
		62082	=>	22114,
		62083	=>	22117,
		62084	=>	22120,
		62085	=>	22123,
		62086	=>	22126,
		62087	=>	22129,
		62088	=>	22132,
		62089	=>	22135,
		62090	=>	22138,
		62091	=>	22141,
		62092	=>	22144,
		62093	=>	22147,
		62094	=>	22149,
		62095	=>	22152,
		62096	=>	22155,
		62097	=>	22158,
		62098	=>	22161,
		62099	=>	22164,
		62100	=>	22167,
		62101	=>	22170,
		62102	=>	22173,
		62103	=>	22176,
		62104	=>	22179,
		62105	=>	22182,
		62106	=>	22185,
		62107	=>	22188,
		62108	=>	22191,
		62109	=>	22194,
		62110	=>	22197,
		62111	=>	22200,
		62112	=>	22203,
		62113	=>	22206,
		62114	=>	22209,
		62115	=>	22212,
		62116	=>	22215,
		62117	=>	22218,
		62118	=>	22221,
		62119	=>	22224,
		62120	=>	22227,
		62121	=>	22230,
		62122	=>	22233,
		62123	=>	22236,
		62124	=>	22239,
		62125	=>	22242,
		62126	=>	22245,
		62127	=>	22248,
		62128	=>	22251,
		62129	=>	22254,
		62130	=>	22257,
		62131	=>	22260,
		62132	=>	22263,
		62133	=>	22265,
		62134	=>	22268,
		62135	=>	22271,
		62136	=>	22274,
		62137	=>	22277,
		62138	=>	22280,
		62139	=>	22283,
		62140	=>	22286,
		62141	=>	22289,
		62142	=>	22292,
		62143	=>	22295,
		62144	=>	22298,
		62145	=>	22301,
		62146	=>	22304,
		62147	=>	22307,
		62148	=>	22310,
		62149	=>	22313,
		62150	=>	22316,
		62151	=>	22319,
		62152	=>	22322,
		62153	=>	22325,
		62154	=>	22328,
		62155	=>	22331,
		62156	=>	22334,
		62157	=>	22337,
		62158	=>	22340,
		62159	=>	22343,
		62160	=>	22346,
		62161	=>	22349,
		62162	=>	22352,
		62163	=>	22355,
		62164	=>	22358,
		62165	=>	22361,
		62166	=>	22364,
		62167	=>	22367,
		62168	=>	22370,
		62169	=>	22373,
		62170	=>	22376,
		62171	=>	22379,
		62172	=>	22382,
		62173	=>	22385,
		62174	=>	22388,
		62175	=>	22391,
		62176	=>	22394,
		62177	=>	22397,
		62178	=>	22399,
		62179	=>	22402,
		62180	=>	22405,
		62181	=>	22408,
		62182	=>	22411,
		62183	=>	22414,
		62184	=>	22417,
		62185	=>	22420,
		62186	=>	22423,
		62187	=>	22426,
		62188	=>	22429,
		62189	=>	22432,
		62190	=>	22435,
		62191	=>	22438,
		62192	=>	22441,
		62193	=>	22444,
		62194	=>	22447,
		62195	=>	22450,
		62196	=>	22453,
		62197	=>	22456,
		62198	=>	22459,
		62199	=>	22462,
		62200	=>	22465,
		62201	=>	22468,
		62202	=>	22471,
		62203	=>	22474,
		62204	=>	22477,
		62205	=>	22480,
		62206	=>	22483,
		62207	=>	22486,
		62208	=>	22489,
		62209	=>	22492,
		62210	=>	22495,
		62211	=>	22498,
		62212	=>	22501,
		62213	=>	22504,
		62214	=>	22507,
		62215	=>	22510,
		62216	=>	22513,
		62217	=>	22516,
		62218	=>	22519,
		62219	=>	22522,
		62220	=>	22525,
		62221	=>	22528,
		62222	=>	22531,
		62223	=>	22534,
		62224	=>	22537,
		62225	=>	22540,
		62226	=>	22543,
		62227	=>	22546,
		62228	=>	22549,
		62229	=>	22552,
		62230	=>	22555,
		62231	=>	22558,
		62232	=>	22561,
		62233	=>	22564,
		62234	=>	22567,
		62235	=>	22570,
		62236	=>	22572,
		62237	=>	22575,
		62238	=>	22578,
		62239	=>	22581,
		62240	=>	22584,
		62241	=>	22587,
		62242	=>	22590,
		62243	=>	22593,
		62244	=>	22596,
		62245	=>	22599,
		62246	=>	22602,
		62247	=>	22605,
		62248	=>	22608,
		62249	=>	22611,
		62250	=>	22614,
		62251	=>	22617,
		62252	=>	22620,
		62253	=>	22623,
		62254	=>	22626,
		62255	=>	22629,
		62256	=>	22632,
		62257	=>	22635,
		62258	=>	22638,
		62259	=>	22641,
		62260	=>	22644,
		62261	=>	22647,
		62262	=>	22650,
		62263	=>	22653,
		62264	=>	22656,
		62265	=>	22659,
		62266	=>	22662,
		62267	=>	22665,
		62268	=>	22668,
		62269	=>	22671,
		62270	=>	22674,
		62271	=>	22677,
		62272	=>	22680,
		62273	=>	22683,
		62274	=>	22686,
		62275	=>	22689,
		62276	=>	22692,
		62277	=>	22695,
		62278	=>	22698,
		62279	=>	22701,
		62280	=>	22704,
		62281	=>	22707,
		62282	=>	22710,
		62283	=>	22713,
		62284	=>	22716,
		62285	=>	22719,
		62286	=>	22722,
		62287	=>	22725,
		62288	=>	22728,
		62289	=>	22731,
		62290	=>	22734,
		62291	=>	22737,
		62292	=>	22740,
		62293	=>	22743,
		62294	=>	22746,
		62295	=>	22749,
		62296	=>	22752,
		62297	=>	22755,
		62298	=>	22758,
		62299	=>	22761,
		62300	=>	22764,
		62301	=>	22767,
		62302	=>	22770,
		62303	=>	22773,
		62304	=>	22776,
		62305	=>	22779,
		62306	=>	22782,
		62307	=>	22785,
		62308	=>	22788,
		62309	=>	22791,
		62310	=>	22794,
		62311	=>	22797,
		62312	=>	22800,
		62313	=>	22803,
		62314	=>	22806,
		62315	=>	22809,
		62316	=>	22812,
		62317	=>	22815,
		62318	=>	22818,
		62319	=>	22821,
		62320	=>	22824,
		62321	=>	22827,
		62322	=>	22830,
		62323	=>	22833,
		62324	=>	22836,
		62325	=>	22839,
		62326	=>	22842,
		62327	=>	22845,
		62328	=>	22848,
		62329	=>	22851,
		62330	=>	22854,
		62331	=>	22857,
		62332	=>	22860,
		62333	=>	22863,
		62334	=>	22866,
		62335	=>	22869,
		62336	=>	22872,
		62337	=>	22875,
		62338	=>	22878,
		62339	=>	22881,
		62340	=>	22884,
		62341	=>	22886,
		62342	=>	22889,
		62343	=>	22892,
		62344	=>	22895,
		62345	=>	22898,
		62346	=>	22901,
		62347	=>	22904,
		62348	=>	22907,
		62349	=>	22910,
		62350	=>	22913,
		62351	=>	22916,
		62352	=>	22919,
		62353	=>	22922,
		62354	=>	22925,
		62355	=>	22928,
		62356	=>	22931,
		62357	=>	22934,
		62358	=>	22937,
		62359	=>	22940,
		62360	=>	22943,
		62361	=>	22946,
		62362	=>	22949,
		62363	=>	22952,
		62364	=>	22955,
		62365	=>	22958,
		62366	=>	22961,
		62367	=>	22964,
		62368	=>	22967,
		62369	=>	22970,
		62370	=>	22973,
		62371	=>	22976,
		62372	=>	22979,
		62373	=>	22982,
		62374	=>	22985,
		62375	=>	22988,
		62376	=>	22991,
		62377	=>	22994,
		62378	=>	22997,
		62379	=>	23000,
		62380	=>	23003,
		62381	=>	23006,
		62382	=>	23009,
		62383	=>	23012,
		62384	=>	23015,
		62385	=>	23018,
		62386	=>	23021,
		62387	=>	23024,
		62388	=>	23027,
		62389	=>	23030,
		62390	=>	23033,
		62391	=>	23036,
		62392	=>	23039,
		62393	=>	23042,
		62394	=>	23045,
		62395	=>	23048,
		62396	=>	23051,
		62397	=>	23054,
		62398	=>	23057,
		62399	=>	23060,
		62400	=>	23063,
		62401	=>	23066,
		62402	=>	23069,
		62403	=>	23072,
		62404	=>	23075,
		62405	=>	23078,
		62406	=>	23081,
		62407	=>	23084,
		62408	=>	23087,
		62409	=>	23090,
		62410	=>	23093,
		62411	=>	23096,
		62412	=>	23099,
		62413	=>	23102,
		62414	=>	23105,
		62415	=>	23108,
		62416	=>	23111,
		62417	=>	23114,
		62418	=>	23117,
		62419	=>	23120,
		62420	=>	23123,
		62421	=>	23126,
		62422	=>	23129,
		62423	=>	23132,
		62424	=>	23135,
		62425	=>	23138,
		62426	=>	23141,
		62427	=>	23144,
		62428	=>	23147,
		62429	=>	23150,
		62430	=>	23153,
		62431	=>	23156,
		62432	=>	23159,
		62433	=>	23162,
		62434	=>	23165,
		62435	=>	23168,
		62436	=>	23171,
		62437	=>	23174,
		62438	=>	23177,
		62439	=>	23180,
		62440	=>	23183,
		62441	=>	23186,
		62442	=>	23189,
		62443	=>	23192,
		62444	=>	23195,
		62445	=>	23198,
		62446	=>	23201,
		62447	=>	23205,
		62448	=>	23208,
		62449	=>	23211,
		62450	=>	23214,
		62451	=>	23217,
		62452	=>	23220,
		62453	=>	23223,
		62454	=>	23226,
		62455	=>	23229,
		62456	=>	23232,
		62457	=>	23235,
		62458	=>	23238,
		62459	=>	23241,
		62460	=>	23244,
		62461	=>	23247,
		62462	=>	23250,
		62463	=>	23253,
		62464	=>	23256,
		62465	=>	23259,
		62466	=>	23262,
		62467	=>	23265,
		62468	=>	23268,
		62469	=>	23271,
		62470	=>	23274,
		62471	=>	23277,
		62472	=>	23280,
		62473	=>	23283,
		62474	=>	23286,
		62475	=>	23289,
		62476	=>	23292,
		62477	=>	23295,
		62478	=>	23298,
		62479	=>	23301,
		62480	=>	23304,
		62481	=>	23307,
		62482	=>	23310,
		62483	=>	23313,
		62484	=>	23316,
		62485	=>	23319,
		62486	=>	23322,
		62487	=>	23325,
		62488	=>	23328,
		62489	=>	23331,
		62490	=>	23334,
		62491	=>	23337,
		62492	=>	23340,
		62493	=>	23343,
		62494	=>	23346,
		62495	=>	23349,
		62496	=>	23352,
		62497	=>	23355,
		62498	=>	23358,
		62499	=>	23361,
		62500	=>	23364,
		62501	=>	23367,
		62502	=>	23370,
		62503	=>	23373,
		62504	=>	23376,
		62505	=>	23379,
		62506	=>	23382,
		62507	=>	23385,
		62508	=>	23388,
		62509	=>	23391,
		62510	=>	23394,
		62511	=>	23397,
		62512	=>	23400,
		62513	=>	23403,
		62514	=>	23406,
		62515	=>	23409,
		62516	=>	23412,
		62517	=>	23415,
		62518	=>	23418,
		62519	=>	23421,
		62520	=>	23424,
		62521	=>	23427,
		62522	=>	23430,
		62523	=>	23433,
		62524	=>	23436,
		62525	=>	23439,
		62526	=>	23442,
		62527	=>	23445,
		62528	=>	23448,
		62529	=>	23451,
		62530	=>	23454,
		62531	=>	23457,
		62532	=>	23460,
		62533	=>	23463,
		62534	=>	23466,
		62535	=>	23469,
		62536	=>	23472,
		62537	=>	23475,
		62538	=>	23478,
		62539	=>	23481,
		62540	=>	23484,
		62541	=>	23487,
		62542	=>	23490,
		62543	=>	23493,
		62544	=>	23496,
		62545	=>	23499,
		62546	=>	23502,
		62547	=>	23505,
		62548	=>	23508,
		62549	=>	23511,
		62550	=>	23514,
		62551	=>	23517,
		62552	=>	23520,
		62553	=>	23523,
		62554	=>	23527,
		62555	=>	23530,
		62556	=>	23533,
		62557	=>	23536,
		62558	=>	23539,
		62559	=>	23542,
		62560	=>	23545,
		62561	=>	23548,
		62562	=>	23551,
		62563	=>	23554,
		62564	=>	23557,
		62565	=>	23560,
		62566	=>	23563,
		62567	=>	23566,
		62568	=>	23569,
		62569	=>	23572,
		62570	=>	23575,
		62571	=>	23578,
		62572	=>	23581,
		62573	=>	23584,
		62574	=>	23587,
		62575	=>	23590,
		62576	=>	23593,
		62577	=>	23596,
		62578	=>	23599,
		62579	=>	23602,
		62580	=>	23605,
		62581	=>	23608,
		62582	=>	23611,
		62583	=>	23614,
		62584	=>	23617,
		62585	=>	23620,
		62586	=>	23623,
		62587	=>	23626,
		62588	=>	23629,
		62589	=>	23632,
		62590	=>	23635,
		62591	=>	23638,
		62592	=>	23641,
		62593	=>	23644,
		62594	=>	23647,
		62595	=>	23650,
		62596	=>	23653,
		62597	=>	23656,
		62598	=>	23659,
		62599	=>	23662,
		62600	=>	23665,
		62601	=>	23668,
		62602	=>	23671,
		62603	=>	23674,
		62604	=>	23677,
		62605	=>	23680,
		62606	=>	23683,
		62607	=>	23686,
		62608	=>	23689,
		62609	=>	23692,
		62610	=>	23695,
		62611	=>	23698,
		62612	=>	23701,
		62613	=>	23704,
		62614	=>	23708,
		62615	=>	23711,
		62616	=>	23714,
		62617	=>	23717,
		62618	=>	23720,
		62619	=>	23723,
		62620	=>	23726,
		62621	=>	23729,
		62622	=>	23732,
		62623	=>	23735,
		62624	=>	23738,
		62625	=>	23741,
		62626	=>	23744,
		62627	=>	23747,
		62628	=>	23750,
		62629	=>	23753,
		62630	=>	23756,
		62631	=>	23759,
		62632	=>	23762,
		62633	=>	23765,
		62634	=>	23768,
		62635	=>	23771,
		62636	=>	23774,
		62637	=>	23777,
		62638	=>	23780,
		62639	=>	23783,
		62640	=>	23786,
		62641	=>	23789,
		62642	=>	23792,
		62643	=>	23795,
		62644	=>	23798,
		62645	=>	23801,
		62646	=>	23804,
		62647	=>	23807,
		62648	=>	23810,
		62649	=>	23813,
		62650	=>	23816,
		62651	=>	23819,
		62652	=>	23822,
		62653	=>	23825,
		62654	=>	23828,
		62655	=>	23831,
		62656	=>	23834,
		62657	=>	23837,
		62658	=>	23840,
		62659	=>	23843,
		62660	=>	23846,
		62661	=>	23849,
		62662	=>	23853,
		62663	=>	23856,
		62664	=>	23859,
		62665	=>	23862,
		62666	=>	23865,
		62667	=>	23868,
		62668	=>	23871,
		62669	=>	23874,
		62670	=>	23877,
		62671	=>	23880,
		62672	=>	23883,
		62673	=>	23886,
		62674	=>	23889,
		62675	=>	23892,
		62676	=>	23895,
		62677	=>	23898,
		62678	=>	23901,
		62679	=>	23904,
		62680	=>	23907,
		62681	=>	23910,
		62682	=>	23913,
		62683	=>	23916,
		62684	=>	23919,
		62685	=>	23922,
		62686	=>	23925,
		62687	=>	23928,
		62688	=>	23931,
		62689	=>	23934,
		62690	=>	23937,
		62691	=>	23940,
		62692	=>	23943,
		62693	=>	23946,
		62694	=>	23949,
		62695	=>	23952,
		62696	=>	23955,
		62697	=>	23958,
		62698	=>	23961,
		62699	=>	23964,
		62700	=>	23967,
		62701	=>	23970,
		62702	=>	23974,
		62703	=>	23977,
		62704	=>	23980,
		62705	=>	23983,
		62706	=>	23986,
		62707	=>	23989,
		62708	=>	23992,
		62709	=>	23995,
		62710	=>	23998,
		62711	=>	24001,
		62712	=>	24004,
		62713	=>	24007,
		62714	=>	24010,
		62715	=>	24013,
		62716	=>	24016,
		62717	=>	24019,
		62718	=>	24022,
		62719	=>	24025,
		62720	=>	24028,
		62721	=>	24031,
		62722	=>	24034,
		62723	=>	24037,
		62724	=>	24040,
		62725	=>	24043,
		62726	=>	24046,
		62727	=>	24049,
		62728	=>	24052,
		62729	=>	24055,
		62730	=>	24058,
		62731	=>	24061,
		62732	=>	24064,
		62733	=>	24067,
		62734	=>	24070,
		62735	=>	24073,
		62736	=>	24076,
		62737	=>	24079,
		62738	=>	24083,
		62739	=>	24086,
		62740	=>	24089,
		62741	=>	24092,
		62742	=>	24095,
		62743	=>	24098,
		62744	=>	24101,
		62745	=>	24104,
		62746	=>	24107,
		62747	=>	24110,
		62748	=>	24113,
		62749	=>	24116,
		62750	=>	24119,
		62751	=>	24122,
		62752	=>	24125,
		62753	=>	24128,
		62754	=>	24131,
		62755	=>	24134,
		62756	=>	24137,
		62757	=>	24140,
		62758	=>	24143,
		62759	=>	24146,
		62760	=>	24149,
		62761	=>	24152,
		62762	=>	24155,
		62763	=>	24158,
		62764	=>	24161,
		62765	=>	24164,
		62766	=>	24167,
		62767	=>	24170,
		62768	=>	24173,
		62769	=>	24176,
		62770	=>	24179,
		62771	=>	24183,
		62772	=>	24186,
		62773	=>	24189,
		62774	=>	24192,
		62775	=>	24195,
		62776	=>	24198,
		62777	=>	24201,
		62778	=>	24204,
		62779	=>	24207,
		62780	=>	24210,
		62781	=>	24213,
		62782	=>	24216,
		62783	=>	24219,
		62784	=>	24222,
		62785	=>	24225,
		62786	=>	24228,
		62787	=>	24231,
		62788	=>	24234,
		62789	=>	24237,
		62790	=>	24240,
		62791	=>	24243,
		62792	=>	24246,
		62793	=>	24249,
		62794	=>	24252,
		62795	=>	24255,
		62796	=>	24258,
		62797	=>	24261,
		62798	=>	24264,
		62799	=>	24267,
		62800	=>	24270,
		62801	=>	24273,
		62802	=>	24277,
		62803	=>	24280,
		62804	=>	24283,
		62805	=>	24286,
		62806	=>	24289,
		62807	=>	24292,
		62808	=>	24295,
		62809	=>	24298,
		62810	=>	24301,
		62811	=>	24304,
		62812	=>	24307,
		62813	=>	24310,
		62814	=>	24313,
		62815	=>	24316,
		62816	=>	24319,
		62817	=>	24322,
		62818	=>	24325,
		62819	=>	24328,
		62820	=>	24331,
		62821	=>	24334,
		62822	=>	24337,
		62823	=>	24340,
		62824	=>	24343,
		62825	=>	24346,
		62826	=>	24349,
		62827	=>	24352,
		62828	=>	24355,
		62829	=>	24358,
		62830	=>	24362,
		62831	=>	24365,
		62832	=>	24368,
		62833	=>	24371,
		62834	=>	24374,
		62835	=>	24377,
		62836	=>	24380,
		62837	=>	24383,
		62838	=>	24386,
		62839	=>	24389,
		62840	=>	24392,
		62841	=>	24395,
		62842	=>	24398,
		62843	=>	24401,
		62844	=>	24404,
		62845	=>	24407,
		62846	=>	24410,
		62847	=>	24413,
		62848	=>	24416,
		62849	=>	24419,
		62850	=>	24422,
		62851	=>	24425,
		62852	=>	24428,
		62853	=>	24431,
		62854	=>	24434,
		62855	=>	24437,
		62856	=>	24440,
		62857	=>	24444,
		62858	=>	24447,
		62859	=>	24450,
		62860	=>	24453,
		62861	=>	24456,
		62862	=>	24459,
		62863	=>	24462,
		62864	=>	24465,
		62865	=>	24468,
		62866	=>	24471,
		62867	=>	24474,
		62868	=>	24477,
		62869	=>	24480,
		62870	=>	24483,
		62871	=>	24486,
		62872	=>	24489,
		62873	=>	24492,
		62874	=>	24495,
		62875	=>	24498,
		62876	=>	24501,
		62877	=>	24504,
		62878	=>	24507,
		62879	=>	24510,
		62880	=>	24513,
		62881	=>	24516,
		62882	=>	24520,
		62883	=>	24523,
		62884	=>	24526,
		62885	=>	24529,
		62886	=>	24532,
		62887	=>	24535,
		62888	=>	24538,
		62889	=>	24541,
		62890	=>	24544,
		62891	=>	24547,
		62892	=>	24550,
		62893	=>	24553,
		62894	=>	24556,
		62895	=>	24559,
		62896	=>	24562,
		62897	=>	24565,
		62898	=>	24568,
		62899	=>	24571,
		62900	=>	24574,
		62901	=>	24577,
		62902	=>	24580,
		62903	=>	24583,
		62904	=>	24586,
		62905	=>	24589,
		62906	=>	24593,
		62907	=>	24596,
		62908	=>	24599,
		62909	=>	24602,
		62910	=>	24605,
		62911	=>	24608,
		62912	=>	24611,
		62913	=>	24614,
		62914	=>	24617,
		62915	=>	24620,
		62916	=>	24623,
		62917	=>	24626,
		62918	=>	24629,
		62919	=>	24632,
		62920	=>	24635,
		62921	=>	24638,
		62922	=>	24641,
		62923	=>	24644,
		62924	=>	24647,
		62925	=>	24650,
		62926	=>	24653,
		62927	=>	24656,
		62928	=>	24659,
		62929	=>	24663,
		62930	=>	24666,
		62931	=>	24669,
		62932	=>	24672,
		62933	=>	24675,
		62934	=>	24678,
		62935	=>	24681,
		62936	=>	24684,
		62937	=>	24687,
		62938	=>	24690,
		62939	=>	24693,
		62940	=>	24696,
		62941	=>	24699,
		62942	=>	24702,
		62943	=>	24705,
		62944	=>	24708,
		62945	=>	24711,
		62946	=>	24714,
		62947	=>	24717,
		62948	=>	24720,
		62949	=>	24723,
		62950	=>	24726,
		62951	=>	24729,
		62952	=>	24733,
		62953	=>	24736,
		62954	=>	24739,
		62955	=>	24742,
		62956	=>	24745,
		62957	=>	24748,
		62958	=>	24751,
		62959	=>	24754,
		62960	=>	24757,
		62961	=>	24760,
		62962	=>	24763,
		62963	=>	24766,
		62964	=>	24769,
		62965	=>	24772,
		62966	=>	24775,
		62967	=>	24778,
		62968	=>	24781,
		62969	=>	24784,
		62970	=>	24787,
		62971	=>	24790,
		62972	=>	24793,
		62973	=>	24797,
		62974	=>	24800,
		62975	=>	24803,
		62976	=>	24806,
		62977	=>	24809,
		62978	=>	24812,
		62979	=>	24815,
		62980	=>	24818,
		62981	=>	24821,
		62982	=>	24824,
		62983	=>	24827,
		62984	=>	24830,
		62985	=>	24833,
		62986	=>	24836,
		62987	=>	24839,
		62988	=>	24842,
		62989	=>	24845,
		62990	=>	24848,
		62991	=>	24851,
		62992	=>	24854,
		62993	=>	24857,
		62994	=>	24861,
		62995	=>	24864,
		62996	=>	24867,
		62997	=>	24870,
		62998	=>	24873,
		62999	=>	24876,
		63000	=>	24879,
		63001	=>	24882,
		63002	=>	24885,
		63003	=>	24888,
		63004	=>	24891,
		63005	=>	24894,
		63006	=>	24897,
		63007	=>	24900,
		63008	=>	24903,
		63009	=>	24906,
		63010	=>	24909,
		63011	=>	24912,
		63012	=>	24915,
		63013	=>	24918,
		63014	=>	24922,
		63015	=>	24925,
		63016	=>	24928,
		63017	=>	24931,
		63018	=>	24934,
		63019	=>	24937,
		63020	=>	24940,
		63021	=>	24943,
		63022	=>	24946,
		63023	=>	24949,
		63024	=>	24952,
		63025	=>	24955,
		63026	=>	24958,
		63027	=>	24961,
		63028	=>	24964,
		63029	=>	24967,
		63030	=>	24970,
		63031	=>	24973,
		63032	=>	24976,
		63033	=>	24979,
		63034	=>	24983,
		63035	=>	24986,
		63036	=>	24989,
		63037	=>	24992,
		63038	=>	24995,
		63039	=>	24998,
		63040	=>	25001,
		63041	=>	25004,
		63042	=>	25007,
		63043	=>	25010,
		63044	=>	25013,
		63045	=>	25016,
		63046	=>	25019,
		63047	=>	25022,
		63048	=>	25025,
		63049	=>	25028,
		63050	=>	25031,
		63051	=>	25034,
		63052	=>	25037,
		63053	=>	25041,
		63054	=>	25044,
		63055	=>	25047,
		63056	=>	25050,
		63057	=>	25053,
		63058	=>	25056,
		63059	=>	25059,
		63060	=>	25062,
		63061	=>	25065,
		63062	=>	25068,
		63063	=>	25071,
		63064	=>	25074,
		63065	=>	25077,
		63066	=>	25080,
		63067	=>	25083,
		63068	=>	25086,
		63069	=>	25089,
		63070	=>	25092,
		63071	=>	25095,
		63072	=>	25099,
		63073	=>	25102,
		63074	=>	25105,
		63075	=>	25108,
		63076	=>	25111,
		63077	=>	25114,
		63078	=>	25117,
		63079	=>	25120,
		63080	=>	25123,
		63081	=>	25126,
		63082	=>	25129,
		63083	=>	25132,
		63084	=>	25135,
		63085	=>	25138,
		63086	=>	25141,
		63087	=>	25144,
		63088	=>	25147,
		63089	=>	25150,
		63090	=>	25154,
		63091	=>	25157,
		63092	=>	25160,
		63093	=>	25163,
		63094	=>	25166,
		63095	=>	25169,
		63096	=>	25172,
		63097	=>	25175,
		63098	=>	25178,
		63099	=>	25181,
		63100	=>	25184,
		63101	=>	25187,
		63102	=>	25190,
		63103	=>	25193,
		63104	=>	25196,
		63105	=>	25199,
		63106	=>	25202,
		63107	=>	25205,
		63108	=>	25209,
		63109	=>	25212,
		63110	=>	25215,
		63111	=>	25218,
		63112	=>	25221,
		63113	=>	25224,
		63114	=>	25227,
		63115	=>	25230,
		63116	=>	25233,
		63117	=>	25236,
		63118	=>	25239,
		63119	=>	25242,
		63120	=>	25245,
		63121	=>	25248,
		63122	=>	25251,
		63123	=>	25254,
		63124	=>	25257,
		63125	=>	25261,
		63126	=>	25264,
		63127	=>	25267,
		63128	=>	25270,
		63129	=>	25273,
		63130	=>	25276,
		63131	=>	25279,
		63132	=>	25282,
		63133	=>	25285,
		63134	=>	25288,
		63135	=>	25291,
		63136	=>	25294,
		63137	=>	25297,
		63138	=>	25300,
		63139	=>	25303,
		63140	=>	25306,
		63141	=>	25309,
		63142	=>	25313,
		63143	=>	25316,
		63144	=>	25319,
		63145	=>	25322,
		63146	=>	25325,
		63147	=>	25328,
		63148	=>	25331,
		63149	=>	25334,
		63150	=>	25337,
		63151	=>	25340,
		63152	=>	25343,
		63153	=>	25346,
		63154	=>	25349,
		63155	=>	25352,
		63156	=>	25355,
		63157	=>	25358,
		63158	=>	25361,
		63159	=>	25365,
		63160	=>	25368,
		63161	=>	25371,
		63162	=>	25374,
		63163	=>	25377,
		63164	=>	25380,
		63165	=>	25383,
		63166	=>	25386,
		63167	=>	25389,
		63168	=>	25392,
		63169	=>	25395,
		63170	=>	25398,
		63171	=>	25401,
		63172	=>	25404,
		63173	=>	25407,
		63174	=>	25410,
		63175	=>	25413,
		63176	=>	25417,
		63177	=>	25420,
		63178	=>	25423,
		63179	=>	25426,
		63180	=>	25429,
		63181	=>	25432,
		63182	=>	25435,
		63183	=>	25438,
		63184	=>	25441,
		63185	=>	25444,
		63186	=>	25447,
		63187	=>	25450,
		63188	=>	25453,
		63189	=>	25456,
		63190	=>	25459,
		63191	=>	25462,
		63192	=>	25466,
		63193	=>	25469,
		63194	=>	25472,
		63195	=>	25475,
		63196	=>	25478,
		63197	=>	25481,
		63198	=>	25484,
		63199	=>	25487,
		63200	=>	25490,
		63201	=>	25493,
		63202	=>	25496,
		63203	=>	25499,
		63204	=>	25502,
		63205	=>	25505,
		63206	=>	25508,
		63207	=>	25511,
		63208	=>	25515,
		63209	=>	25518,
		63210	=>	25521,
		63211	=>	25524,
		63212	=>	25527,
		63213	=>	25530,
		63214	=>	25533,
		63215	=>	25536,
		63216	=>	25539,
		63217	=>	25542,
		63218	=>	25545,
		63219	=>	25548,
		63220	=>	25551,
		63221	=>	25554,
		63222	=>	25557,
		63223	=>	25561,
		63224	=>	25564,
		63225	=>	25567,
		63226	=>	25570,
		63227	=>	25573,
		63228	=>	25576,
		63229	=>	25579,
		63230	=>	25582,
		63231	=>	25585,
		63232	=>	25588,
		63233	=>	25591,
		63234	=>	25594,
		63235	=>	25597,
		63236	=>	25600,
		63237	=>	25603,
		63238	=>	25606,
		63239	=>	25610,
		63240	=>	25613,
		63241	=>	25616,
		63242	=>	25619,
		63243	=>	25622,
		63244	=>	25625,
		63245	=>	25628,
		63246	=>	25631,
		63247	=>	25634,
		63248	=>	25637,
		63249	=>	25640,
		63250	=>	25643,
		63251	=>	25646,
		63252	=>	25649,
		63253	=>	25652,
		63254	=>	25656,
		63255	=>	25659,
		63256	=>	25662,
		63257	=>	25665,
		63258	=>	25668,
		63259	=>	25671,
		63260	=>	25674,
		63261	=>	25677,
		63262	=>	25680,
		63263	=>	25683,
		63264	=>	25686,
		63265	=>	25689,
		63266	=>	25692,
		63267	=>	25695,
		63268	=>	25698,
		63269	=>	25702,
		63270	=>	25705,
		63271	=>	25708,
		63272	=>	25711,
		63273	=>	25714,
		63274	=>	25717,
		63275	=>	25720,
		63276	=>	25723,
		63277	=>	25726,
		63278	=>	25729,
		63279	=>	25732,
		63280	=>	25735,
		63281	=>	25738,
		63282	=>	25741,
		63283	=>	25745,
		63284	=>	25748,
		63285	=>	25751,
		63286	=>	25754,
		63287	=>	25757,
		63288	=>	25760,
		63289	=>	25763,
		63290	=>	25766,
		63291	=>	25769,
		63292	=>	25772,
		63293	=>	25775,
		63294	=>	25778,
		63295	=>	25781,
		63296	=>	25784,
		63297	=>	25787,
		63298	=>	25791,
		63299	=>	25794,
		63300	=>	25797,
		63301	=>	25800,
		63302	=>	25803,
		63303	=>	25806,
		63304	=>	25809,
		63305	=>	25812,
		63306	=>	25815,
		63307	=>	25818,
		63308	=>	25821,
		63309	=>	25824,
		63310	=>	25827,
		63311	=>	25830,
		63312	=>	25834,
		63313	=>	25837,
		63314	=>	25840,
		63315	=>	25843,
		63316	=>	25846,
		63317	=>	25849,
		63318	=>	25852,
		63319	=>	25855,
		63320	=>	25858,
		63321	=>	25861,
		63322	=>	25864,
		63323	=>	25867,
		63324	=>	25870,
		63325	=>	25873,
		63326	=>	25877,
		63327	=>	25880,
		63328	=>	25883,
		63329	=>	25886,
		63330	=>	25889,
		63331	=>	25892,
		63332	=>	25895,
		63333	=>	25898,
		63334	=>	25901,
		63335	=>	25904,
		63336	=>	25907,
		63337	=>	25910,
		63338	=>	25913,
		63339	=>	25916,
		63340	=>	25920,
		63341	=>	25923,
		63342	=>	25926,
		63343	=>	25929,
		63344	=>	25932,
		63345	=>	25935,
		63346	=>	25938,
		63347	=>	25941,
		63348	=>	25944,
		63349	=>	25947,
		63350	=>	25950,
		63351	=>	25953,
		63352	=>	25956,
		63353	=>	25959,
		63354	=>	25963,
		63355	=>	25966,
		63356	=>	25969,
		63357	=>	25972,
		63358	=>	25975,
		63359	=>	25978,
		63360	=>	25981,
		63361	=>	25984,
		63362	=>	25987,
		63363	=>	25990,
		63364	=>	25993,
		63365	=>	25996,
		63366	=>	25999,
		63367	=>	26002,
		63368	=>	26006,
		63369	=>	26009,
		63370	=>	26012,
		63371	=>	26015,
		63372	=>	26018,
		63373	=>	26021,
		63374	=>	26024,
		63375	=>	26027,
		63376	=>	26030,
		63377	=>	26033,
		63378	=>	26036,
		63379	=>	26039,
		63380	=>	26042,
		63381	=>	26046,
		63382	=>	26049,
		63383	=>	26052,
		63384	=>	26055,
		63385	=>	26058,
		63386	=>	26061,
		63387	=>	26064,
		63388	=>	26067,
		63389	=>	26070,
		63390	=>	26073,
		63391	=>	26076,
		63392	=>	26079,
		63393	=>	26082,
		63394	=>	26086,
		63395	=>	26089,
		63396	=>	26092,
		63397	=>	26095,
		63398	=>	26098,
		63399	=>	26101,
		63400	=>	26104,
		63401	=>	26107,
		63402	=>	26110,
		63403	=>	26113,
		63404	=>	26116,
		63405	=>	26119,
		63406	=>	26122,
		63407	=>	26125,
		63408	=>	26129,
		63409	=>	26132,
		63410	=>	26135,
		63411	=>	26138,
		63412	=>	26141,
		63413	=>	26144,
		63414	=>	26147,
		63415	=>	26150,
		63416	=>	26153,
		63417	=>	26156,
		63418	=>	26159,
		63419	=>	26162,
		63420	=>	26165,
		63421	=>	26169,
		63422	=>	26172,
		63423	=>	26175,
		63424	=>	26178,
		63425	=>	26181,
		63426	=>	26184,
		63427	=>	26187,
		63428	=>	26190,
		63429	=>	26193,
		63430	=>	26196,
		63431	=>	26199,
		63432	=>	26202,
		63433	=>	26206,
		63434	=>	26209,
		63435	=>	26212,
		63436	=>	26215,
		63437	=>	26218,
		63438	=>	26221,
		63439	=>	26224,
		63440	=>	26227,
		63441	=>	26230,
		63442	=>	26233,
		63443	=>	26236,
		63444	=>	26239,
		63445	=>	26242,
		63446	=>	26246,
		63447	=>	26249,
		63448	=>	26252,
		63449	=>	26255,
		63450	=>	26258,
		63451	=>	26261,
		63452	=>	26264,
		63453	=>	26267,
		63454	=>	26270,
		63455	=>	26273,
		63456	=>	26276,
		63457	=>	26279,
		63458	=>	26282,
		63459	=>	26286,
		63460	=>	26289,
		63461	=>	26292,
		63462	=>	26295,
		63463	=>	26298,
		63464	=>	26301,
		63465	=>	26304,
		63466	=>	26307,
		63467	=>	26310,
		63468	=>	26313,
		63469	=>	26316,
		63470	=>	26319,
		63471	=>	26323,
		63472	=>	26326,
		63473	=>	26329,
		63474	=>	26332,
		63475	=>	26335,
		63476	=>	26338,
		63477	=>	26341,
		63478	=>	26344,
		63479	=>	26347,
		63480	=>	26350,
		63481	=>	26353,
		63482	=>	26356,
		63483	=>	26359,
		63484	=>	26363,
		63485	=>	26366,
		63486	=>	26369,
		63487	=>	26372,
		63488	=>	26375,
		63489	=>	26378,
		63490	=>	26381,
		63491	=>	26384,
		63492	=>	26387,
		63493	=>	26390,
		63494	=>	26393,
		63495	=>	26396,
		63496	=>	26400,
		63497	=>	26403,
		63498	=>	26406,
		63499	=>	26409,
		63500	=>	26412,
		63501	=>	26415,
		63502	=>	26418,
		63503	=>	26421,
		63504	=>	26424,
		63505	=>	26427,
		63506	=>	26430,
		63507	=>	26433,
		63508	=>	26437,
		63509	=>	26440,
		63510	=>	26443,
		63511	=>	26446,
		63512	=>	26449,
		63513	=>	26452,
		63514	=>	26455,
		63515	=>	26458,
		63516	=>	26461,
		63517	=>	26464,
		63518	=>	26467,
		63519	=>	26470,
		63520	=>	26474,
		63521	=>	26477,
		63522	=>	26480,
		63523	=>	26483,
		63524	=>	26486,
		63525	=>	26489,
		63526	=>	26492,
		63527	=>	26495,
		63528	=>	26498,
		63529	=>	26501,
		63530	=>	26504,
		63531	=>	26507,
		63532	=>	26511,
		63533	=>	26514,
		63534	=>	26517,
		63535	=>	26520,
		63536	=>	26523,
		63537	=>	26526,
		63538	=>	26529,
		63539	=>	26532,
		63540	=>	26535,
		63541	=>	26538,
		63542	=>	26541,
		63543	=>	26544,
		63544	=>	26548,
		63545	=>	26551,
		63546	=>	26554,
		63547	=>	26557,
		63548	=>	26560,
		63549	=>	26563,
		63550	=>	26566,
		63551	=>	26569,
		63552	=>	26572,
		63553	=>	26575,
		63554	=>	26578,
		63555	=>	26581,
		63556	=>	26585,
		63557	=>	26588,
		63558	=>	26591,
		63559	=>	26594,
		63560	=>	26597,
		63561	=>	26600,
		63562	=>	26603,
		63563	=>	26606,
		63564	=>	26609,
		63565	=>	26612,
		63566	=>	26615,
		63567	=>	26618,
		63568	=>	26622,
		63569	=>	26625,
		63570	=>	26628,
		63571	=>	26631,
		63572	=>	26634,
		63573	=>	26637,
		63574	=>	26640,
		63575	=>	26643,
		63576	=>	26646,
		63577	=>	26649,
		63578	=>	26652,
		63579	=>	26656,
		63580	=>	26659,
		63581	=>	26662,
		63582	=>	26665,
		63583	=>	26668,
		63584	=>	26671,
		63585	=>	26674,
		63586	=>	26677,
		63587	=>	26680,
		63588	=>	26683,
		63589	=>	26686,
		63590	=>	26689,
		63591	=>	26693,
		63592	=>	26696,
		63593	=>	26699,
		63594	=>	26702,
		63595	=>	26705,
		63596	=>	26708,
		63597	=>	26711,
		63598	=>	26714,
		63599	=>	26717,
		63600	=>	26720,
		63601	=>	26723,
		63602	=>	26727,
		63603	=>	26730,
		63604	=>	26733,
		63605	=>	26736,
		63606	=>	26739,
		63607	=>	26742,
		63608	=>	26745,
		63609	=>	26748,
		63610	=>	26751,
		63611	=>	26754,
		63612	=>	26757,
		63613	=>	26760,
		63614	=>	26764,
		63615	=>	26767,
		63616	=>	26770,
		63617	=>	26773,
		63618	=>	26776,
		63619	=>	26779,
		63620	=>	26782,
		63621	=>	26785,
		63622	=>	26788,
		63623	=>	26791,
		63624	=>	26794,
		63625	=>	26798,
		63626	=>	26801,
		63627	=>	26804,
		63628	=>	26807,
		63629	=>	26810,
		63630	=>	26813,
		63631	=>	26816,
		63632	=>	26819,
		63633	=>	26822,
		63634	=>	26825,
		63635	=>	26828,
		63636	=>	26832,
		63637	=>	26835,
		63638	=>	26838,
		63639	=>	26841,
		63640	=>	26844,
		63641	=>	26847,
		63642	=>	26850,
		63643	=>	26853,
		63644	=>	26856,
		63645	=>	26859,
		63646	=>	26862,
		63647	=>	26866,
		63648	=>	26869,
		63649	=>	26872,
		63650	=>	26875,
		63651	=>	26878,
		63652	=>	26881,
		63653	=>	26884,
		63654	=>	26887,
		63655	=>	26890,
		63656	=>	26893,
		63657	=>	26896,
		63658	=>	26900,
		63659	=>	26903,
		63660	=>	26906,
		63661	=>	26909,
		63662	=>	26912,
		63663	=>	26915,
		63664	=>	26918,
		63665	=>	26921,
		63666	=>	26924,
		63667	=>	26927,
		63668	=>	26930,
		63669	=>	26934,
		63670	=>	26937,
		63671	=>	26940,
		63672	=>	26943,
		63673	=>	26946,
		63674	=>	26949,
		63675	=>	26952,
		63676	=>	26955,
		63677	=>	26958,
		63678	=>	26961,
		63679	=>	26964,
		63680	=>	26968,
		63681	=>	26971,
		63682	=>	26974,
		63683	=>	26977,
		63684	=>	26980,
		63685	=>	26983,
		63686	=>	26986,
		63687	=>	26989,
		63688	=>	26992,
		63689	=>	26995,
		63690	=>	26998,
		63691	=>	27002,
		63692	=>	27005,
		63693	=>	27008,
		63694	=>	27011,
		63695	=>	27014,
		63696	=>	27017,
		63697	=>	27020,
		63698	=>	27023,
		63699	=>	27026,
		63700	=>	27029,
		63701	=>	27032,
		63702	=>	27036,
		63703	=>	27039,
		63704	=>	27042,
		63705	=>	27045,
		63706	=>	27048,
		63707	=>	27051,
		63708	=>	27054,
		63709	=>	27057,
		63710	=>	27060,
		63711	=>	27063,
		63712	=>	27066,
		63713	=>	27070,
		63714	=>	27073,
		63715	=>	27076,
		63716	=>	27079,
		63717	=>	27082,
		63718	=>	27085,
		63719	=>	27088,
		63720	=>	27091,
		63721	=>	27094,
		63722	=>	27097,
		63723	=>	27101,
		63724	=>	27104,
		63725	=>	27107,
		63726	=>	27110,
		63727	=>	27113,
		63728	=>	27116,
		63729	=>	27119,
		63730	=>	27122,
		63731	=>	27125,
		63732	=>	27128,
		63733	=>	27131,
		63734	=>	27135,
		63735	=>	27138,
		63736	=>	27141,
		63737	=>	27144,
		63738	=>	27147,
		63739	=>	27150,
		63740	=>	27153,
		63741	=>	27156,
		63742	=>	27159,
		63743	=>	27162,
		63744	=>	27166,
		63745	=>	27169,
		63746	=>	27172,
		63747	=>	27175,
		63748	=>	27178,
		63749	=>	27181,
		63750	=>	27184,
		63751	=>	27187,
		63752	=>	27190,
		63753	=>	27193,
		63754	=>	27196,
		63755	=>	27200,
		63756	=>	27203,
		63757	=>	27206,
		63758	=>	27209,
		63759	=>	27212,
		63760	=>	27215,
		63761	=>	27218,
		63762	=>	27221,
		63763	=>	27224,
		63764	=>	27227,
		63765	=>	27231,
		63766	=>	27234,
		63767	=>	27237,
		63768	=>	27240,
		63769	=>	27243,
		63770	=>	27246,
		63771	=>	27249,
		63772	=>	27252,
		63773	=>	27255,
		63774	=>	27258,
		63775	=>	27261,
		63776	=>	27265,
		63777	=>	27268,
		63778	=>	27271,
		63779	=>	27274,
		63780	=>	27277,
		63781	=>	27280,
		63782	=>	27283,
		63783	=>	27286,
		63784	=>	27289,
		63785	=>	27292,
		63786	=>	27296,
		63787	=>	27299,
		63788	=>	27302,
		63789	=>	27305,
		63790	=>	27308,
		63791	=>	27311,
		63792	=>	27314,
		63793	=>	27317,
		63794	=>	27320,
		63795	=>	27323,
		63796	=>	27327,
		63797	=>	27330,
		63798	=>	27333,
		63799	=>	27336,
		63800	=>	27339,
		63801	=>	27342,
		63802	=>	27345,
		63803	=>	27348,
		63804	=>	27351,
		63805	=>	27354,
		63806	=>	27358,
		63807	=>	27361,
		63808	=>	27364,
		63809	=>	27367,
		63810	=>	27370,
		63811	=>	27373,
		63812	=>	27376,
		63813	=>	27379,
		63814	=>	27382,
		63815	=>	27385,
		63816	=>	27388,
		63817	=>	27392,
		63818	=>	27395,
		63819	=>	27398,
		63820	=>	27401,
		63821	=>	27404,
		63822	=>	27407,
		63823	=>	27410,
		63824	=>	27413,
		63825	=>	27416,
		63826	=>	27419,
		63827	=>	27423,
		63828	=>	27426,
		63829	=>	27429,
		63830	=>	27432,
		63831	=>	27435,
		63832	=>	27438,
		63833	=>	27441,
		63834	=>	27444,
		63835	=>	27447,
		63836	=>	27450,
		63837	=>	27454,
		63838	=>	27457,
		63839	=>	27460,
		63840	=>	27463,
		63841	=>	27466,
		63842	=>	27469,
		63843	=>	27472,
		63844	=>	27475,
		63845	=>	27478,
		63846	=>	27481,
		63847	=>	27485,
		63848	=>	27488,
		63849	=>	27491,
		63850	=>	27494,
		63851	=>	27497,
		63852	=>	27500,
		63853	=>	27503,
		63854	=>	27506,
		63855	=>	27509,
		63856	=>	27512,
		63857	=>	27516,
		63858	=>	27519,
		63859	=>	27522,
		63860	=>	27525,
		63861	=>	27528,
		63862	=>	27531,
		63863	=>	27534,
		63864	=>	27537,
		63865	=>	27540,
		63866	=>	27544,
		63867	=>	27547,
		63868	=>	27550,
		63869	=>	27553,
		63870	=>	27556,
		63871	=>	27559,
		63872	=>	27562,
		63873	=>	27565,
		63874	=>	27568,
		63875	=>	27571,
		63876	=>	27575,
		63877	=>	27578,
		63878	=>	27581,
		63879	=>	27584,
		63880	=>	27587,
		63881	=>	27590,
		63882	=>	27593,
		63883	=>	27596,
		63884	=>	27599,
		63885	=>	27602,
		63886	=>	27606,
		63887	=>	27609,
		63888	=>	27612,
		63889	=>	27615,
		63890	=>	27618,
		63891	=>	27621,
		63892	=>	27624,
		63893	=>	27627,
		63894	=>	27630,
		63895	=>	27633,
		63896	=>	27637,
		63897	=>	27640,
		63898	=>	27643,
		63899	=>	27646,
		63900	=>	27649,
		63901	=>	27652,
		63902	=>	27655,
		63903	=>	27658,
		63904	=>	27661,
		63905	=>	27664,
		63906	=>	27668,
		63907	=>	27671,
		63908	=>	27674,
		63909	=>	27677,
		63910	=>	27680,
		63911	=>	27683,
		63912	=>	27686,
		63913	=>	27689,
		63914	=>	27692,
		63915	=>	27696,
		63916	=>	27699,
		63917	=>	27702,
		63918	=>	27705,
		63919	=>	27708,
		63920	=>	27711,
		63921	=>	27714,
		63922	=>	27717,
		63923	=>	27720,
		63924	=>	27723,
		63925	=>	27727,
		63926	=>	27730,
		63927	=>	27733,
		63928	=>	27736,
		63929	=>	27739,
		63930	=>	27742,
		63931	=>	27745,
		63932	=>	27748,
		63933	=>	27751,
		63934	=>	27755,
		63935	=>	27758,
		63936	=>	27761,
		63937	=>	27764,
		63938	=>	27767,
		63939	=>	27770,
		63940	=>	27773,
		63941	=>	27776,
		63942	=>	27779,
		63943	=>	27782,
		63944	=>	27786,
		63945	=>	27789,
		63946	=>	27792,
		63947	=>	27795,
		63948	=>	27798,
		63949	=>	27801,
		63950	=>	27804,
		63951	=>	27807,
		63952	=>	27810,
		63953	=>	27814,
		63954	=>	27817,
		63955	=>	27820,
		63956	=>	27823,
		63957	=>	27826,
		63958	=>	27829,
		63959	=>	27832,
		63960	=>	27835,
		63961	=>	27838,
		63962	=>	27841,
		63963	=>	27845,
		63964	=>	27848,
		63965	=>	27851,
		63966	=>	27854,
		63967	=>	27857,
		63968	=>	27860,
		63969	=>	27863,
		63970	=>	27866,
		63971	=>	27869,
		63972	=>	27873,
		63973	=>	27876,
		63974	=>	27879,
		63975	=>	27882,
		63976	=>	27885,
		63977	=>	27888,
		63978	=>	27891,
		63979	=>	27894,
		63980	=>	27897,
		63981	=>	27900,
		63982	=>	27904,
		63983	=>	27907,
		63984	=>	27910,
		63985	=>	27913,
		63986	=>	27916,
		63987	=>	27919,
		63988	=>	27922,
		63989	=>	27925,
		63990	=>	27928,
		63991	=>	27932,
		63992	=>	27935,
		63993	=>	27938,
		63994	=>	27941,
		63995	=>	27944,
		63996	=>	27947,
		63997	=>	27950,
		63998	=>	27953,
		63999	=>	27956,
		64000	=>	27960,
		64001	=>	27963,
		64002	=>	27966,
		64003	=>	27969,
		64004	=>	27972,
		64005	=>	27975,
		64006	=>	27978,
		64007	=>	27981,
		64008	=>	27984,
		64009	=>	27987,
		64010	=>	27991,
		64011	=>	27994,
		64012	=>	27997,
		64013	=>	28000,
		64014	=>	28003,
		64015	=>	28006,
		64016	=>	28009,
		64017	=>	28012,
		64018	=>	28015,
		64019	=>	28019,
		64020	=>	28022,
		64021	=>	28025,
		64022	=>	28028,
		64023	=>	28031,
		64024	=>	28034,
		64025	=>	28037,
		64026	=>	28040,
		64027	=>	28043,
		64028	=>	28047,
		64029	=>	28050,
		64030	=>	28053,
		64031	=>	28056,
		64032	=>	28059,
		64033	=>	28062,
		64034	=>	28065,
		64035	=>	28068,
		64036	=>	28071,
		64037	=>	28075,
		64038	=>	28078,
		64039	=>	28081,
		64040	=>	28084,
		64041	=>	28087,
		64042	=>	28090,
		64043	=>	28093,
		64044	=>	28096,
		64045	=>	28099,
		64046	=>	28103,
		64047	=>	28106,
		64048	=>	28109,
		64049	=>	28112,
		64050	=>	28115,
		64051	=>	28118,
		64052	=>	28121,
		64053	=>	28124,
		64054	=>	28127,
		64055	=>	28130,
		64056	=>	28134,
		64057	=>	28137,
		64058	=>	28140,
		64059	=>	28143,
		64060	=>	28146,
		64061	=>	28149,
		64062	=>	28152,
		64063	=>	28155,
		64064	=>	28158,
		64065	=>	28162,
		64066	=>	28165,
		64067	=>	28168,
		64068	=>	28171,
		64069	=>	28174,
		64070	=>	28177,
		64071	=>	28180,
		64072	=>	28183,
		64073	=>	28186,
		64074	=>	28190,
		64075	=>	28193,
		64076	=>	28196,
		64077	=>	28199,
		64078	=>	28202,
		64079	=>	28205,
		64080	=>	28208,
		64081	=>	28211,
		64082	=>	28214,
		64083	=>	28218,
		64084	=>	28221,
		64085	=>	28224,
		64086	=>	28227,
		64087	=>	28230,
		64088	=>	28233,
		64089	=>	28236,
		64090	=>	28239,
		64091	=>	28242,
		64092	=>	28246,
		64093	=>	28249,
		64094	=>	28252,
		64095	=>	28255,
		64096	=>	28258,
		64097	=>	28261,
		64098	=>	28264,
		64099	=>	28267,
		64100	=>	28270,
		64101	=>	28274,
		64102	=>	28277,
		64103	=>	28280,
		64104	=>	28283,
		64105	=>	28286,
		64106	=>	28289,
		64107	=>	28292,
		64108	=>	28295,
		64109	=>	28298,
		64110	=>	28302,
		64111	=>	28305,
		64112	=>	28308,
		64113	=>	28311,
		64114	=>	28314,
		64115	=>	28317,
		64116	=>	28320,
		64117	=>	28323,
		64118	=>	28326,
		64119	=>	28330,
		64120	=>	28333,
		64121	=>	28336,
		64122	=>	28339,
		64123	=>	28342,
		64124	=>	28345,
		64125	=>	28348,
		64126	=>	28351,
		64127	=>	28355,
		64128	=>	28358,
		64129	=>	28361,
		64130	=>	28364,
		64131	=>	28367,
		64132	=>	28370,
		64133	=>	28373,
		64134	=>	28376,
		64135	=>	28379,
		64136	=>	28383,
		64137	=>	28386,
		64138	=>	28389,
		64139	=>	28392,
		64140	=>	28395,
		64141	=>	28398,
		64142	=>	28401,
		64143	=>	28404,
		64144	=>	28407,
		64145	=>	28411,
		64146	=>	28414,
		64147	=>	28417,
		64148	=>	28420,
		64149	=>	28423,
		64150	=>	28426,
		64151	=>	28429,
		64152	=>	28432,
		64153	=>	28435,
		64154	=>	28439,
		64155	=>	28442,
		64156	=>	28445,
		64157	=>	28448,
		64158	=>	28451,
		64159	=>	28454,
		64160	=>	28457,
		64161	=>	28460,
		64162	=>	28463,
		64163	=>	28467,
		64164	=>	28470,
		64165	=>	28473,
		64166	=>	28476,
		64167	=>	28479,
		64168	=>	28482,
		64169	=>	28485,
		64170	=>	28488,
		64171	=>	28492,
		64172	=>	28495,
		64173	=>	28498,
		64174	=>	28501,
		64175	=>	28504,
		64176	=>	28507,
		64177	=>	28510,
		64178	=>	28513,
		64179	=>	28516,
		64180	=>	28520,
		64181	=>	28523,
		64182	=>	28526,
		64183	=>	28529,
		64184	=>	28532,
		64185	=>	28535,
		64186	=>	28538,
		64187	=>	28541,
		64188	=>	28544,
		64189	=>	28548,
		64190	=>	28551,
		64191	=>	28554,
		64192	=>	28557,
		64193	=>	28560,
		64194	=>	28563,
		64195	=>	28566,
		64196	=>	28569,
		64197	=>	28573,
		64198	=>	28576,
		64199	=>	28579,
		64200	=>	28582,
		64201	=>	28585,
		64202	=>	28588,
		64203	=>	28591,
		64204	=>	28594,
		64205	=>	28597,
		64206	=>	28601,
		64207	=>	28604,
		64208	=>	28607,
		64209	=>	28610,
		64210	=>	28613,
		64211	=>	28616,
		64212	=>	28619,
		64213	=>	28622,
		64214	=>	28625,
		64215	=>	28629,
		64216	=>	28632,
		64217	=>	28635,
		64218	=>	28638,
		64219	=>	28641,
		64220	=>	28644,
		64221	=>	28647,
		64222	=>	28650,
		64223	=>	28654,
		64224	=>	28657,
		64225	=>	28660,
		64226	=>	28663,
		64227	=>	28666,
		64228	=>	28669,
		64229	=>	28672,
		64230	=>	28675,
		64231	=>	28678,
		64232	=>	28682,
		64233	=>	28685,
		64234	=>	28688,
		64235	=>	28691,
		64236	=>	28694,
		64237	=>	28697,
		64238	=>	28700,
		64239	=>	28703,
		64240	=>	28707,
		64241	=>	28710,
		64242	=>	28713,
		64243	=>	28716,
		64244	=>	28719,
		64245	=>	28722,
		64246	=>	28725,
		64247	=>	28728,
		64248	=>	28731,
		64249	=>	28735,
		64250	=>	28738,
		64251	=>	28741,
		64252	=>	28744,
		64253	=>	28747,
		64254	=>	28750,
		64255	=>	28753,
		64256	=>	28756,
		64257	=>	28760,
		64258	=>	28763,
		64259	=>	28766,
		64260	=>	28769,
		64261	=>	28772,
		64262	=>	28775,
		64263	=>	28778,
		64264	=>	28781,
		64265	=>	28784,
		64266	=>	28788,
		64267	=>	28791,
		64268	=>	28794,
		64269	=>	28797,
		64270	=>	28800,
		64271	=>	28803,
		64272	=>	28806,
		64273	=>	28809,
		64274	=>	28813,
		64275	=>	28816,
		64276	=>	28819,
		64277	=>	28822,
		64278	=>	28825,
		64279	=>	28828,
		64280	=>	28831,
		64281	=>	28834,
		64282	=>	28837,
		64283	=>	28841,
		64284	=>	28844,
		64285	=>	28847,
		64286	=>	28850,
		64287	=>	28853,
		64288	=>	28856,
		64289	=>	28859,
		64290	=>	28862,
		64291	=>	28866,
		64292	=>	28869,
		64293	=>	28872,
		64294	=>	28875,
		64295	=>	28878,
		64296	=>	28881,
		64297	=>	28884,
		64298	=>	28887,
		64299	=>	28891,
		64300	=>	28894,
		64301	=>	28897,
		64302	=>	28900,
		64303	=>	28903,
		64304	=>	28906,
		64305	=>	28909,
		64306	=>	28912,
		64307	=>	28915,
		64308	=>	28919,
		64309	=>	28922,
		64310	=>	28925,
		64311	=>	28928,
		64312	=>	28931,
		64313	=>	28934,
		64314	=>	28937,
		64315	=>	28940,
		64316	=>	28944,
		64317	=>	28947,
		64318	=>	28950,
		64319	=>	28953,
		64320	=>	28956,
		64321	=>	28959,
		64322	=>	28962,
		64323	=>	28965,
		64324	=>	28969,
		64325	=>	28972,
		64326	=>	28975,
		64327	=>	28978,
		64328	=>	28981,
		64329	=>	28984,
		64330	=>	28987,
		64331	=>	28990,
		64332	=>	28993,
		64333	=>	28997,
		64334	=>	29000,
		64335	=>	29003,
		64336	=>	29006,
		64337	=>	29009,
		64338	=>	29012,
		64339	=>	29015,
		64340	=>	29018,
		64341	=>	29022,
		64342	=>	29025,
		64343	=>	29028,
		64344	=>	29031,
		64345	=>	29034,
		64346	=>	29037,
		64347	=>	29040,
		64348	=>	29043,
		64349	=>	29047,
		64350	=>	29050,
		64351	=>	29053,
		64352	=>	29056,
		64353	=>	29059,
		64354	=>	29062,
		64355	=>	29065,
		64356	=>	29068,
		64357	=>	29072,
		64358	=>	29075,
		64359	=>	29078,
		64360	=>	29081,
		64361	=>	29084,
		64362	=>	29087,
		64363	=>	29090,
		64364	=>	29093,
		64365	=>	29096,
		64366	=>	29100,
		64367	=>	29103,
		64368	=>	29106,
		64369	=>	29109,
		64370	=>	29112,
		64371	=>	29115,
		64372	=>	29118,
		64373	=>	29121,
		64374	=>	29125,
		64375	=>	29128,
		64376	=>	29131,
		64377	=>	29134,
		64378	=>	29137,
		64379	=>	29140,
		64380	=>	29143,
		64381	=>	29146,
		64382	=>	29150,
		64383	=>	29153,
		64384	=>	29156,
		64385	=>	29159,
		64386	=>	29162,
		64387	=>	29165,
		64388	=>	29168,
		64389	=>	29171,
		64390	=>	29175,
		64391	=>	29178,
		64392	=>	29181,
		64393	=>	29184,
		64394	=>	29187,
		64395	=>	29190,
		64396	=>	29193,
		64397	=>	29196,
		64398	=>	29200,
		64399	=>	29203,
		64400	=>	29206,
		64401	=>	29209,
		64402	=>	29212,
		64403	=>	29215,
		64404	=>	29218,
		64405	=>	29221,
		64406	=>	29224,
		64407	=>	29228,
		64408	=>	29231,
		64409	=>	29234,
		64410	=>	29237,
		64411	=>	29240,
		64412	=>	29243,
		64413	=>	29246,
		64414	=>	29249,
		64415	=>	29253,
		64416	=>	29256,
		64417	=>	29259,
		64418	=>	29262,
		64419	=>	29265,
		64420	=>	29268,
		64421	=>	29271,
		64422	=>	29274,
		64423	=>	29278,
		64424	=>	29281,
		64425	=>	29284,
		64426	=>	29287,
		64427	=>	29290,
		64428	=>	29293,
		64429	=>	29296,
		64430	=>	29299,
		64431	=>	29303,
		64432	=>	29306,
		64433	=>	29309,
		64434	=>	29312,
		64435	=>	29315,
		64436	=>	29318,
		64437	=>	29321,
		64438	=>	29324,
		64439	=>	29328,
		64440	=>	29331,
		64441	=>	29334,
		64442	=>	29337,
		64443	=>	29340,
		64444	=>	29343,
		64445	=>	29346,
		64446	=>	29349,
		64447	=>	29353,
		64448	=>	29356,
		64449	=>	29359,
		64450	=>	29362,
		64451	=>	29365,
		64452	=>	29368,
		64453	=>	29371,
		64454	=>	29374,
		64455	=>	29378,
		64456	=>	29381,
		64457	=>	29384,
		64458	=>	29387,
		64459	=>	29390,
		64460	=>	29393,
		64461	=>	29396,
		64462	=>	29399,
		64463	=>	29403,
		64464	=>	29406,
		64465	=>	29409,
		64466	=>	29412,
		64467	=>	29415,
		64468	=>	29418,
		64469	=>	29421,
		64470	=>	29424,
		64471	=>	29428,
		64472	=>	29431,
		64473	=>	29434,
		64474	=>	29437,
		64475	=>	29440,
		64476	=>	29443,
		64477	=>	29446,
		64478	=>	29449,
		64479	=>	29453,
		64480	=>	29456,
		64481	=>	29459,
		64482	=>	29462,
		64483	=>	29465,
		64484	=>	29468,
		64485	=>	29471,
		64486	=>	29474,
		64487	=>	29478,
		64488	=>	29481,
		64489	=>	29484,
		64490	=>	29487,
		64491	=>	29490,
		64492	=>	29493,
		64493	=>	29496,
		64494	=>	29499,
		64495	=>	29503,
		64496	=>	29506,
		64497	=>	29509,
		64498	=>	29512,
		64499	=>	29515,
		64500	=>	29518,
		64501	=>	29521,
		64502	=>	29524,
		64503	=>	29528,
		64504	=>	29531,
		64505	=>	29534,
		64506	=>	29537,
		64507	=>	29540,
		64508	=>	29543,
		64509	=>	29546,
		64510	=>	29549,
		64511	=>	29553,
		64512	=>	29556,
		64513	=>	29559,
		64514	=>	29562,
		64515	=>	29565,
		64516	=>	29568,
		64517	=>	29571,
		64518	=>	29574,
		64519	=>	29578,
		64520	=>	29581,
		64521	=>	29584,
		64522	=>	29587,
		64523	=>	29590,
		64524	=>	29593,
		64525	=>	29596,
		64526	=>	29599,
		64527	=>	29603,
		64528	=>	29606,
		64529	=>	29609,
		64530	=>	29612,
		64531	=>	29615,
		64532	=>	29618,
		64533	=>	29621,
		64534	=>	29625,
		64535	=>	29628,
		64536	=>	29631,
		64537	=>	29634,
		64538	=>	29637,
		64539	=>	29640,
		64540	=>	29643,
		64541	=>	29646,
		64542	=>	29650,
		64543	=>	29653,
		64544	=>	29656,
		64545	=>	29659,
		64546	=>	29662,
		64547	=>	29665,
		64548	=>	29668,
		64549	=>	29671,
		64550	=>	29675,
		64551	=>	29678,
		64552	=>	29681,
		64553	=>	29684,
		64554	=>	29687,
		64555	=>	29690,
		64556	=>	29693,
		64557	=>	29696,
		64558	=>	29700,
		64559	=>	29703,
		64560	=>	29706,
		64561	=>	29709,
		64562	=>	29712,
		64563	=>	29715,
		64564	=>	29718,
		64565	=>	29721,
		64566	=>	29725,
		64567	=>	29728,
		64568	=>	29731,
		64569	=>	29734,
		64570	=>	29737,
		64571	=>	29740,
		64572	=>	29743,
		64573	=>	29746,
		64574	=>	29750,
		64575	=>	29753,
		64576	=>	29756,
		64577	=>	29759,
		64578	=>	29762,
		64579	=>	29765,
		64580	=>	29768,
		64581	=>	29772,
		64582	=>	29775,
		64583	=>	29778,
		64584	=>	29781,
		64585	=>	29784,
		64586	=>	29787,
		64587	=>	29790,
		64588	=>	29793,
		64589	=>	29797,
		64590	=>	29800,
		64591	=>	29803,
		64592	=>	29806,
		64593	=>	29809,
		64594	=>	29812,
		64595	=>	29815,
		64596	=>	29818,
		64597	=>	29822,
		64598	=>	29825,
		64599	=>	29828,
		64600	=>	29831,
		64601	=>	29834,
		64602	=>	29837,
		64603	=>	29840,
		64604	=>	29843,
		64605	=>	29847,
		64606	=>	29850,
		64607	=>	29853,
		64608	=>	29856,
		64609	=>	29859,
		64610	=>	29862,
		64611	=>	29865,
		64612	=>	29869,
		64613	=>	29872,
		64614	=>	29875,
		64615	=>	29878,
		64616	=>	29881,
		64617	=>	29884,
		64618	=>	29887,
		64619	=>	29890,
		64620	=>	29894,
		64621	=>	29897,
		64622	=>	29900,
		64623	=>	29903,
		64624	=>	29906,
		64625	=>	29909,
		64626	=>	29912,
		64627	=>	29915,
		64628	=>	29919,
		64629	=>	29922,
		64630	=>	29925,
		64631	=>	29928,
		64632	=>	29931,
		64633	=>	29934,
		64634	=>	29937,
		64635	=>	29940,
		64636	=>	29944,
		64637	=>	29947,
		64638	=>	29950,
		64639	=>	29953,
		64640	=>	29956,
		64641	=>	29959,
		64642	=>	29962,
		64643	=>	29966,
		64644	=>	29969,
		64645	=>	29972,
		64646	=>	29975,
		64647	=>	29978,
		64648	=>	29981,
		64649	=>	29984,
		64650	=>	29987,
		64651	=>	29991,
		64652	=>	29994,
		64653	=>	29997,
		64654	=>	30000,
		64655	=>	30003,
		64656	=>	30006,
		64657	=>	30009,
		64658	=>	30012,
		64659	=>	30016,
		64660	=>	30019,
		64661	=>	30022,
		64662	=>	30025,
		64663	=>	30028,
		64664	=>	30031,
		64665	=>	30034,
		64666	=>	30038,
		64667	=>	30041,
		64668	=>	30044,
		64669	=>	30047,
		64670	=>	30050,
		64671	=>	30053,
		64672	=>	30056,
		64673	=>	30059,
		64674	=>	30063,
		64675	=>	30066,
		64676	=>	30069,
		64677	=>	30072,
		64678	=>	30075,
		64679	=>	30078,
		64680	=>	30081,
		64681	=>	30084,
		64682	=>	30088,
		64683	=>	30091,
		64684	=>	30094,
		64685	=>	30097,
		64686	=>	30100,
		64687	=>	30103,
		64688	=>	30106,
		64689	=>	30110,
		64690	=>	30113,
		64691	=>	30116,
		64692	=>	30119,
		64693	=>	30122,
		64694	=>	30125,
		64695	=>	30128,
		64696	=>	30131,
		64697	=>	30135,
		64698	=>	30138,
		64699	=>	30141,
		64700	=>	30144,
		64701	=>	30147,
		64702	=>	30150,
		64703	=>	30153,
		64704	=>	30157,
		64705	=>	30160,
		64706	=>	30163,
		64707	=>	30166,
		64708	=>	30169,
		64709	=>	30172,
		64710	=>	30175,
		64711	=>	30178,
		64712	=>	30182,
		64713	=>	30185,
		64714	=>	30188,
		64715	=>	30191,
		64716	=>	30194,
		64717	=>	30197,
		64718	=>	30200,
		64719	=>	30203,
		64720	=>	30207,
		64721	=>	30210,
		64722	=>	30213,
		64723	=>	30216,
		64724	=>	30219,
		64725	=>	30222,
		64726	=>	30225,
		64727	=>	30229,
		64728	=>	30232,
		64729	=>	30235,
		64730	=>	30238,
		64731	=>	30241,
		64732	=>	30244,
		64733	=>	30247,
		64734	=>	30250,
		64735	=>	30254,
		64736	=>	30257,
		64737	=>	30260,
		64738	=>	30263,
		64739	=>	30266,
		64740	=>	30269,
		64741	=>	30272,
		64742	=>	30276,
		64743	=>	30279,
		64744	=>	30282,
		64745	=>	30285,
		64746	=>	30288,
		64747	=>	30291,
		64748	=>	30294,
		64749	=>	30297,
		64750	=>	30301,
		64751	=>	30304,
		64752	=>	30307,
		64753	=>	30310,
		64754	=>	30313,
		64755	=>	30316,
		64756	=>	30319,
		64757	=>	30323,
		64758	=>	30326,
		64759	=>	30329,
		64760	=>	30332,
		64761	=>	30335,
		64762	=>	30338,
		64763	=>	30341,
		64764	=>	30344,
		64765	=>	30348,
		64766	=>	30351,
		64767	=>	30354,
		64768	=>	30357,
		64769	=>	30360,
		64770	=>	30363,
		64771	=>	30366,
		64772	=>	30370,
		64773	=>	30373,
		64774	=>	30376,
		64775	=>	30379,
		64776	=>	30382,
		64777	=>	30385,
		64778	=>	30388,
		64779	=>	30391,
		64780	=>	30395,
		64781	=>	30398,
		64782	=>	30401,
		64783	=>	30404,
		64784	=>	30407,
		64785	=>	30410,
		64786	=>	30413,
		64787	=>	30417,
		64788	=>	30420,
		64789	=>	30423,
		64790	=>	30426,
		64791	=>	30429,
		64792	=>	30432,
		64793	=>	30435,
		64794	=>	30438,
		64795	=>	30442,
		64796	=>	30445,
		64797	=>	30448,
		64798	=>	30451,
		64799	=>	30454,
		64800	=>	30457,
		64801	=>	30460,
		64802	=>	30464,
		64803	=>	30467,
		64804	=>	30470,
		64805	=>	30473,
		64806	=>	30476,
		64807	=>	30479,
		64808	=>	30482,
		64809	=>	30485,
		64810	=>	30489,
		64811	=>	30492,
		64812	=>	30495,
		64813	=>	30498,
		64814	=>	30501,
		64815	=>	30504,
		64816	=>	30507,
		64817	=>	30511,
		64818	=>	30514,
		64819	=>	30517,
		64820	=>	30520,
		64821	=>	30523,
		64822	=>	30526,
		64823	=>	30529,
		64824	=>	30532,
		64825	=>	30536,
		64826	=>	30539,
		64827	=>	30542,
		64828	=>	30545,
		64829	=>	30548,
		64830	=>	30551,
		64831	=>	30554,
		64832	=>	30558,
		64833	=>	30561,
		64834	=>	30564,
		64835	=>	30567,
		64836	=>	30570,
		64837	=>	30573,
		64838	=>	30576,
		64839	=>	30579,
		64840	=>	30583,
		64841	=>	30586,
		64842	=>	30589,
		64843	=>	30592,
		64844	=>	30595,
		64845	=>	30598,
		64846	=>	30601,
		64847	=>	30605,
		64848	=>	30608,
		64849	=>	30611,
		64850	=>	30614,
		64851	=>	30617,
		64852	=>	30620,
		64853	=>	30623,
		64854	=>	30626,
		64855	=>	30630,
		64856	=>	30633,
		64857	=>	30636,
		64858	=>	30639,
		64859	=>	30642,
		64860	=>	30645,
		64861	=>	30648,
		64862	=>	30652,
		64863	=>	30655,
		64864	=>	30658,
		64865	=>	30661,
		64866	=>	30664,
		64867	=>	30667,
		64868	=>	30670,
		64869	=>	30674,
		64870	=>	30677,
		64871	=>	30680,
		64872	=>	30683,
		64873	=>	30686,
		64874	=>	30689,
		64875	=>	30692,
		64876	=>	30695,
		64877	=>	30699,
		64878	=>	30702,
		64879	=>	30705,
		64880	=>	30708,
		64881	=>	30711,
		64882	=>	30714,
		64883	=>	30717,
		64884	=>	30721,
		64885	=>	30724,
		64886	=>	30727,
		64887	=>	30730,
		64888	=>	30733,
		64889	=>	30736,
		64890	=>	30739,
		64891	=>	30742,
		64892	=>	30746,
		64893	=>	30749,
		64894	=>	30752,
		64895	=>	30755,
		64896	=>	30758,
		64897	=>	30761,
		64898	=>	30764,
		64899	=>	30768,
		64900	=>	30771,
		64901	=>	30774,
		64902	=>	30777,
		64903	=>	30780,
		64904	=>	30783,
		64905	=>	30786,
		64906	=>	30790,
		64907	=>	30793,
		64908	=>	30796,
		64909	=>	30799,
		64910	=>	30802,
		64911	=>	30805,
		64912	=>	30808,
		64913	=>	30811,
		64914	=>	30815,
		64915	=>	30818,
		64916	=>	30821,
		64917	=>	30824,
		64918	=>	30827,
		64919	=>	30830,
		64920	=>	30833,
		64921	=>	30837,
		64922	=>	30840,
		64923	=>	30843,
		64924	=>	30846,
		64925	=>	30849,
		64926	=>	30852,
		64927	=>	30855,
		64928	=>	30859,
		64929	=>	30862,
		64930	=>	30865,
		64931	=>	30868,
		64932	=>	30871,
		64933	=>	30874,
		64934	=>	30877,
		64935	=>	30880,
		64936	=>	30884,
		64937	=>	30887,
		64938	=>	30890,
		64939	=>	30893,
		64940	=>	30896,
		64941	=>	30899,
		64942	=>	30902,
		64943	=>	30906,
		64944	=>	30909,
		64945	=>	30912,
		64946	=>	30915,
		64947	=>	30918,
		64948	=>	30921,
		64949	=>	30924,
		64950	=>	30928,
		64951	=>	30931,
		64952	=>	30934,
		64953	=>	30937,
		64954	=>	30940,
		64955	=>	30943,
		64956	=>	30946,
		64957	=>	30949,
		64958	=>	30953,
		64959	=>	30956,
		64960	=>	30959,
		64961	=>	30962,
		64962	=>	30965,
		64963	=>	30968,
		64964	=>	30971,
		64965	=>	30975,
		64966	=>	30978,
		64967	=>	30981,
		64968	=>	30984,
		64969	=>	30987,
		64970	=>	30990,
		64971	=>	30993,
		64972	=>	30997,
		64973	=>	31000,
		64974	=>	31003,
		64975	=>	31006,
		64976	=>	31009,
		64977	=>	31012,
		64978	=>	31015,
		64979	=>	31018,
		64980	=>	31022,
		64981	=>	31025,
		64982	=>	31028,
		64983	=>	31031,
		64984	=>	31034,
		64985	=>	31037,
		64986	=>	31040,
		64987	=>	31044,
		64988	=>	31047,
		64989	=>	31050,
		64990	=>	31053,
		64991	=>	31056,
		64992	=>	31059,
		64993	=>	31062,
		64994	=>	31066,
		64995	=>	31069,
		64996	=>	31072,
		64997	=>	31075,
		64998	=>	31078,
		64999	=>	31081,
		65000	=>	31084,
		65001	=>	31088,
		65002	=>	31091,
		65003	=>	31094,
		65004	=>	31097,
		65005	=>	31100,
		65006	=>	31103,
		65007	=>	31106,
		65008	=>	31109,
		65009	=>	31113,
		65010	=>	31116,
		65011	=>	31119,
		65012	=>	31122,
		65013	=>	31125,
		65014	=>	31128,
		65015	=>	31131,
		65016	=>	31135,
		65017	=>	31138,
		65018	=>	31141,
		65019	=>	31144,
		65020	=>	31147,
		65021	=>	31150,
		65022	=>	31153,
		65023	=>	31157,
		65024	=>	31160,
		65025	=>	31163,
		65026	=>	31166,
		65027	=>	31169,
		65028	=>	31172,
		65029	=>	31175,
		65030	=>	31179,
		65031	=>	31182,
		65032	=>	31185,
		65033	=>	31188,
		65034	=>	31191,
		65035	=>	31194,
		65036	=>	31197,
		65037	=>	31200,
		65038	=>	31204,
		65039	=>	31207,
		65040	=>	31210,
		65041	=>	31213,
		65042	=>	31216,
		65043	=>	31219,
		65044	=>	31222,
		65045	=>	31226,
		65046	=>	31229,
		65047	=>	31232,
		65048	=>	31235,
		65049	=>	31238,
		65050	=>	31241,
		65051	=>	31244,
		65052	=>	31248,
		65053	=>	31251,
		65054	=>	31254,
		65055	=>	31257,
		65056	=>	31260,
		65057	=>	31263,
		65058	=>	31266,
		65059	=>	31270,
		65060	=>	31273,
		65061	=>	31276,
		65062	=>	31279,
		65063	=>	31282,
		65064	=>	31285,
		65065	=>	31288,
		65066	=>	31291,
		65067	=>	31295,
		65068	=>	31298,
		65069	=>	31301,
		65070	=>	31304,
		65071	=>	31307,
		65072	=>	31310,
		65073	=>	31313,
		65074	=>	31317,
		65075	=>	31320,
		65076	=>	31323,
		65077	=>	31326,
		65078	=>	31329,
		65079	=>	31332,
		65080	=>	31335,
		65081	=>	31339,
		65082	=>	31342,
		65083	=>	31345,
		65084	=>	31348,
		65085	=>	31351,
		65086	=>	31354,
		65087	=>	31357,
		65088	=>	31361,
		65089	=>	31364,
		65090	=>	31367,
		65091	=>	31370,
		65092	=>	31373,
		65093	=>	31376,
		65094	=>	31379,
		65095	=>	31382,
		65096	=>	31386,
		65097	=>	31389,
		65098	=>	31392,
		65099	=>	31395,
		65100	=>	31398,
		65101	=>	31401,
		65102	=>	31404,
		65103	=>	31408,
		65104	=>	31411,
		65105	=>	31414,
		65106	=>	31417,
		65107	=>	31420,
		65108	=>	31423,
		65109	=>	31426,
		65110	=>	31430,
		65111	=>	31433,
		65112	=>	31436,
		65113	=>	31439,
		65114	=>	31442,
		65115	=>	31445,
		65116	=>	31448,
		65117	=>	31452,
		65118	=>	31455,
		65119	=>	31458,
		65120	=>	31461,
		65121	=>	31464,
		65122	=>	31467,
		65123	=>	31470,
		65124	=>	31474,
		65125	=>	31477,
		65126	=>	31480,
		65127	=>	31483,
		65128	=>	31486,
		65129	=>	31489,
		65130	=>	31492,
		65131	=>	31495,
		65132	=>	31499,
		65133	=>	31502,
		65134	=>	31505,
		65135	=>	31508,
		65136	=>	31511,
		65137	=>	31514,
		65138	=>	31517,
		65139	=>	31521,
		65140	=>	31524,
		65141	=>	31527,
		65142	=>	31530,
		65143	=>	31533,
		65144	=>	31536,
		65145	=>	31539,
		65146	=>	31543,
		65147	=>	31546,
		65148	=>	31549,
		65149	=>	31552,
		65150	=>	31555,
		65151	=>	31558,
		65152	=>	31561,
		65153	=>	31565,
		65154	=>	31568,
		65155	=>	31571,
		65156	=>	31574,
		65157	=>	31577,
		65158	=>	31580,
		65159	=>	31583,
		65160	=>	31587,
		65161	=>	31590,
		65162	=>	31593,
		65163	=>	31596,
		65164	=>	31599,
		65165	=>	31602,
		65166	=>	31605,
		65167	=>	31609,
		65168	=>	31612,
		65169	=>	31615,
		65170	=>	31618,
		65171	=>	31621,
		65172	=>	31624,
		65173	=>	31627,
		65174	=>	31630,
		65175	=>	31634,
		65176	=>	31637,
		65177	=>	31640,
		65178	=>	31643,
		65179	=>	31646,
		65180	=>	31649,
		65181	=>	31652,
		65182	=>	31656,
		65183	=>	31659,
		65184	=>	31662,
		65185	=>	31665,
		65186	=>	31668,
		65187	=>	31671,
		65188	=>	31674,
		65189	=>	31678,
		65190	=>	31681,
		65191	=>	31684,
		65192	=>	31687,
		65193	=>	31690,
		65194	=>	31693,
		65195	=>	31696,
		65196	=>	31700,
		65197	=>	31703,
		65198	=>	31706,
		65199	=>	31709,
		65200	=>	31712,
		65201	=>	31715,
		65202	=>	31718,
		65203	=>	31722,
		65204	=>	31725,
		65205	=>	31728,
		65206	=>	31731,
		65207	=>	31734,
		65208	=>	31737,
		65209	=>	31740,
		65210	=>	31744,
		65211	=>	31747,
		65212	=>	31750,
		65213	=>	31753,
		65214	=>	31756,
		65215	=>	31759,
		65216	=>	31762,
		65217	=>	31766,
		65218	=>	31769,
		65219	=>	31772,
		65220	=>	31775,
		65221	=>	31778,
		65222	=>	31781,
		65223	=>	31784,
		65224	=>	31787,
		65225	=>	31791,
		65226	=>	31794,
		65227	=>	31797,
		65228	=>	31800,
		65229	=>	31803,
		65230	=>	31806,
		65231	=>	31809,
		65232	=>	31813,
		65233	=>	31816,
		65234	=>	31819,
		65235	=>	31822,
		65236	=>	31825,
		65237	=>	31828,
		65238	=>	31831,
		65239	=>	31835,
		65240	=>	31838,
		65241	=>	31841,
		65242	=>	31844,
		65243	=>	31847,
		65244	=>	31850,
		65245	=>	31853,
		65246	=>	31857,
		65247	=>	31860,
		65248	=>	31863,
		65249	=>	31866,
		65250	=>	31869,
		65251	=>	31872,
		65252	=>	31875,
		65253	=>	31879,
		65254	=>	31882,
		65255	=>	31885,
		65256	=>	31888,
		65257	=>	31891,
		65258	=>	31894,
		65259	=>	31897,
		65260	=>	31901,
		65261	=>	31904,
		65262	=>	31907,
		65263	=>	31910,
		65264	=>	31913,
		65265	=>	31916,
		65266	=>	31919,
		65267	=>	31923,
		65268	=>	31926,
		65269	=>	31929,
		65270	=>	31932,
		65271	=>	31935,
		65272	=>	31938,
		65273	=>	31941,
		65274	=>	31945,
		65275	=>	31948,
		65276	=>	31951,
		65277	=>	31954,
		65278	=>	31957,
		65279	=>	31960,
		65280	=>	31963,
		65281	=>	31966,
		65282	=>	31970,
		65283	=>	31973,
		65284	=>	31976,
		65285	=>	31979,
		65286	=>	31982,
		65287	=>	31985,
		65288	=>	31988,
		65289	=>	31992,
		65290	=>	31995,
		65291	=>	31998,
		65292	=>	32001,
		65293	=>	32004,
		65294	=>	32007,
		65295	=>	32010,
		65296	=>	32014,
		65297	=>	32017,
		65298	=>	32020,
		65299	=>	32023,
		65300	=>	32026,
		65301	=>	32029,
		65302	=>	32032,
		65303	=>	32036,
		65304	=>	32039,
		65305	=>	32042,
		65306	=>	32045,
		65307	=>	32048,
		65308	=>	32051,
		65309	=>	32054,
		65310	=>	32058,
		65311	=>	32061,
		65312	=>	32064,
		65313	=>	32067,
		65314	=>	32070,
		65315	=>	32073,
		65316	=>	32076,
		65317	=>	32080,
		65318	=>	32083,
		65319	=>	32086,
		65320	=>	32089,
		65321	=>	32092,
		65322	=>	32095,
		65323	=>	32098,
		65324	=>	32102,
		65325	=>	32105,
		65326	=>	32108,
		65327	=>	32111,
		65328	=>	32114,
		65329	=>	32117,
		65330	=>	32120,
		65331	=>	32124,
		65332	=>	32127,
		65333	=>	32130,
		65334	=>	32133,
		65335	=>	32136,
		65336	=>	32139,
		65337	=>	32142,
		65338	=>	32146,
		65339	=>	32149,
		65340	=>	32152,
		65341	=>	32155,
		65342	=>	32158,
		65343	=>	32161,
		65344	=>	32164,
		65345	=>	32167,
		65346	=>	32171,
		65347	=>	32174,
		65348	=>	32177,
		65349	=>	32180,
		65350	=>	32183,
		65351	=>	32186,
		65352	=>	32189,
		65353	=>	32193,
		65354	=>	32196,
		65355	=>	32199,
		65356	=>	32202,
		65357	=>	32205,
		65358	=>	32208,
		65359	=>	32211,
		65360	=>	32215,
		65361	=>	32218,
		65362	=>	32221,
		65363	=>	32224,
		65364	=>	32227,
		65365	=>	32230,
		65366	=>	32233,
		65367	=>	32237,
		65368	=>	32240,
		65369	=>	32243,
		65370	=>	32246,
		65371	=>	32249,
		65372	=>	32252,
		65373	=>	32255,
		65374	=>	32259,
		65375	=>	32262,
		65376	=>	32265,
		65377	=>	32268,
		65378	=>	32271,
		65379	=>	32274,
		65380	=>	32277,
		65381	=>	32281,
		65382	=>	32284,
		65383	=>	32287,
		65384	=>	32290,
		65385	=>	32293,
		65386	=>	32296,
		65387	=>	32299,
		65388	=>	32303,
		65389	=>	32306,
		65390	=>	32309,
		65391	=>	32312,
		65392	=>	32315,
		65393	=>	32318,
		65394	=>	32321,
		65395	=>	32325,
		65396	=>	32328,
		65397	=>	32331,
		65398	=>	32334,
		65399	=>	32337,
		65400	=>	32340,
		65401	=>	32343,
		65402	=>	32347,
		65403	=>	32350,
		65404	=>	32353,
		65405	=>	32356,
		65406	=>	32359,
		65407	=>	32362,
		65408	=>	32365,
		65409	=>	32369,
		65410	=>	32372,
		65411	=>	32375,
		65412	=>	32378,
		65413	=>	32381,
		65414	=>	32384,
		65415	=>	32387,
		65416	=>	32391,
		65417	=>	32394,
		65418	=>	32397,
		65419	=>	32400,
		65420	=>	32403,
		65421	=>	32406,
		65422	=>	32409,
		65423	=>	32413,
		65424	=>	32416,
		65425	=>	32419,
		65426	=>	32422,
		65427	=>	32425,
		65428	=>	32428,
		65429	=>	32431,
		65430	=>	32435,
		65431	=>	32438,
		65432	=>	32441,
		65433	=>	32444,
		65434	=>	32447,
		65435	=>	32450,
		65436	=>	32453,
		65437	=>	32456,
		65438	=>	32460,
		65439	=>	32463,
		65440	=>	32466,
		65441	=>	32469,
		65442	=>	32472,
		65443	=>	32475,
		65444	=>	32478,
		65445	=>	32482,
		65446	=>	32485,
		65447	=>	32488,
		65448	=>	32491,
		65449	=>	32494,
		65450	=>	32497,
		65451	=>	32500,
		65452	=>	32504,
		65453	=>	32507,
		65454	=>	32510,
		65455	=>	32513,
		65456	=>	32516,
		65457	=>	32519,
		65458	=>	32522,
		65459	=>	32526,
		65460	=>	32529,
		65461	=>	32532,
		65462	=>	32535,
		65463	=>	32538,
		65464	=>	32541,
		65465	=>	32544,
		65466	=>	32548,
		65467	=>	32551,
		65468	=>	32554,
		65469	=>	32557,
		65470	=>	32560,
		65471	=>	32563,
		65472	=>	32566,
		65473	=>	32570,
		65474	=>	32573,
		65475	=>	32576,
		65476	=>	32579,
		65477	=>	32582,
		65478	=>	32585,
		65479	=>	32588,
		65480	=>	32592,
		65481	=>	32595,
		65482	=>	32598,
		65483	=>	32601,
		65484	=>	32604,
		65485	=>	32607,
		65486	=>	32610,
		65487	=>	32614,
		65488	=>	32617,
		65489	=>	32620,
		65490	=>	32623,
		65491	=>	32626,
		65492	=>	32629,
		65493	=>	32632,
		65494	=>	32636,
		65495	=>	32639,
		65496	=>	32642,
		65497	=>	32645,
		65498	=>	32648,
		65499	=>	32651,
		65500	=>	32654,
		65501	=>	32658,
		65502	=>	32661,
		65503	=>	32664,
		65504	=>	32667,
		65505	=>	32670,
		65506	=>	32673,
		65507	=>	32676,
		65508	=>	32680,
		65509	=>	32683,
		65510	=>	32686,
		65511	=>	32689,
		65512	=>	32692,
		65513	=>	32695,
		65514	=>	32698,
		65515	=>	32702,
		65516	=>	32705,
		65517	=>	32708,
		65518	=>	32711,
		65519	=>	32714,
		65520	=>	32717,
		65521	=>	32720,
		65522	=>	32724,
		65523	=>	32727,
		65524	=>	32730,
		65525	=>	32733,
		65526	=>	32736,
		65527	=>	32739,
		65528	=>	32742,
		65529	=>	32746,
		65530	=>	32749,
		65531	=>	32752,
		65532	=>	32755,
		65533	=>	32758,
		65534	=>	32761,
		65535	=>	32764

);

begin
	LUT_data <= std_logic_vector(TO_UNSIGNED(LUT(TO_INTEGER(unsigned(LUT_line))), 16));
end rtl;
